--Tabla de consulta de datos
library IEEE;
use IEEE.std_logic_1164.all;

entity LUT_SIN_SIGNAL is
port (
    F	:	in std_logic_vector(11 downto 0);
    s	: 	out std_logic_vector(11 downto 0)
    );
  end LUT_SIN_SIGNAL;
  
  architecture tabla of LUT_SIN_SIGNAL is
 begin
  process(F)
  begin case F is
  when "000000000000"=> s <="100000000000"; -- Argumento 0 Funcion 0.00000000
  when "000000000001"=> s <="100000000011"; -- Argumento 1 Funcion 0.00153398
  when "000000000010"=> s <="100000000110"; -- Argumento 2 Funcion 0.00306796
  when "000000000011"=> s <="100000001001"; -- Argumento 3 Funcion 0.00460193
  when "000000000100"=> s <="100000001100"; -- Argumento 4 Funcion 0.00613588
  when "000000000101"=> s <="100000001111"; -- Argumento 5 Funcion 0.00766983
  when "000000000110"=> s <="100000010010"; -- Argumento 6 Funcion 0.00920375
  when "000000000111"=> s <="100000010101"; -- Argumento 7 Funcion 0.01073766
  when "000000001000"=> s <="100000011001"; -- Argumento 8 Funcion 0.01227154
  when "000000001001"=> s <="100000011100"; -- Argumento 9 Funcion 0.01380539
  when "000000001010"=> s <="100000011111"; -- Argumento 10 Funcion 0.01533921
  when "000000001011"=> s <="100000100010"; -- Argumento 11 Funcion 0.01687299
  when "000000001100"=> s <="100000100101"; -- Argumento 12 Funcion 0.01840673
  when "000000001101"=> s <="100000101000"; -- Argumento 13 Funcion 0.01994043
  when "000000001110"=> s <="100000101011"; -- Argumento 14 Funcion 0.02147408
  when "000000001111"=> s <="100000101111"; -- Argumento 15 Funcion 0.02300768
  when "000000010000"=> s <="100000110010"; -- Argumento 16 Funcion 0.02454123
  when "000000010001"=> s <="100000110101"; -- Argumento 17 Funcion 0.02607472
  when "000000010010"=> s <="100000111000"; -- Argumento 18 Funcion 0.02760815
  when "000000010011"=> s <="100000111011"; -- Argumento 19 Funcion 0.02914151
  when "000000010100"=> s <="100000111110"; -- Argumento 20 Funcion 0.03067480
  when "000000010101"=> s <="100001000001"; -- Argumento 21 Funcion 0.03220803
  when "000000010110"=> s <="100001000101"; -- Argumento 22 Funcion 0.03374117
  when "000000010111"=> s <="100001001000"; -- Argumento 23 Funcion 0.03527424
  when "000000011000"=> s <="100001001011"; -- Argumento 24 Funcion 0.03680722
  when "000000011001"=> s <="100001001110"; -- Argumento 25 Funcion 0.03834012
  when "000000011010"=> s <="100001010001"; -- Argumento 26 Funcion 0.03987293
  when "000000011011"=> s <="100001010100"; -- Argumento 27 Funcion 0.04140564
  when "000000011100"=> s <="100001010111"; -- Argumento 28 Funcion 0.04293826
  when "000000011101"=> s <="100001011011"; -- Argumento 29 Funcion 0.04447077
  when "000000011110"=> s <="100001011110"; -- Argumento 30 Funcion 0.04600318
  when "000000011111"=> s <="100001100001"; -- Argumento 31 Funcion 0.04753548
  when "000000100000"=> s <="100001100100"; -- Argumento 32 Funcion 0.04906767
  when "000000100001"=> s <="100001100111"; -- Argumento 33 Funcion 0.05059975
  when "000000100010"=> s <="100001101010"; -- Argumento 34 Funcion 0.05213170
  when "000000100011"=> s <="100001101101"; -- Argumento 35 Funcion 0.05366354
  when "000000100100"=> s <="100001110001"; -- Argumento 36 Funcion 0.05519524
  when "000000100101"=> s <="100001110100"; -- Argumento 37 Funcion 0.05672682
  when "000000100110"=> s <="100001110111"; -- Argumento 38 Funcion 0.05825826
  when "000000100111"=> s <="100001111010"; -- Argumento 39 Funcion 0.05978957
  when "000000101000"=> s <="100001111101"; -- Argumento 40 Funcion 0.06132074
  when "000000101001"=> s <="100010000000"; -- Argumento 41 Funcion 0.06285176
  when "000000101010"=> s <="100010000011"; -- Argumento 42 Funcion 0.06438263
  when "000000101011"=> s <="100010000110"; -- Argumento 43 Funcion 0.06591335
  when "000000101100"=> s <="100010001010"; -- Argumento 44 Funcion 0.06744392
  when "000000101101"=> s <="100010001101"; -- Argumento 45 Funcion 0.06897433
  when "000000101110"=> s <="100010010000"; -- Argumento 46 Funcion 0.07050457
  when "000000101111"=> s <="100010010011"; -- Argumento 47 Funcion 0.07203465
  when "000000110000"=> s <="100010010110"; -- Argumento 48 Funcion 0.07356456
  when "000000110001"=> s <="100010011001"; -- Argumento 49 Funcion 0.07509430
  when "000000110010"=> s <="100010011100"; -- Argumento 50 Funcion 0.07662386
  when "000000110011"=> s <="100010100000"; -- Argumento 51 Funcion 0.07815324
  when "000000110100"=> s <="100010100011"; -- Argumento 52 Funcion 0.07968244
  when "000000110101"=> s <="100010100110"; -- Argumento 53 Funcion 0.08121145
  when "000000110110"=> s <="100010101001"; -- Argumento 54 Funcion 0.08274026
  when "000000110111"=> s <="100010101100"; -- Argumento 55 Funcion 0.08426889
  when "000000111000"=> s <="100010101111"; -- Argumento 56 Funcion 0.08579731
  when "000000111001"=> s <="100010110010"; -- Argumento 57 Funcion 0.08732554
  when "000000111010"=> s <="100010110101"; -- Argumento 58 Funcion 0.08885355
  when "000000111011"=> s <="100010111001"; -- Argumento 59 Funcion 0.09038136
  when "000000111100"=> s <="100010111100"; -- Argumento 60 Funcion 0.09190896
  when "000000111101"=> s <="100010111111"; -- Argumento 61 Funcion 0.09343634
  when "000000111110"=> s <="100011000010"; -- Argumento 62 Funcion 0.09496350
  when "000000111111"=> s <="100011000101"; -- Argumento 63 Funcion 0.09649043
  when "000001000000"=> s <="100011001000"; -- Argumento 64 Funcion 0.09801714
  when "000001000001"=> s <="100011001011"; -- Argumento 65 Funcion 0.09954362
  when "000001000010"=> s <="100011001110"; -- Argumento 66 Funcion 0.10106986
  when "000001000011"=> s <="100011010010"; -- Argumento 67 Funcion 0.10259587
  when "000001000100"=> s <="100011010101"; -- Argumento 68 Funcion 0.10412163
  when "000001000101"=> s <="100011011000"; -- Argumento 69 Funcion 0.10564715
  when "000001000110"=> s <="100011011011"; -- Argumento 70 Funcion 0.10717242
  when "000001000111"=> s <="100011011110"; -- Argumento 71 Funcion 0.10869744
  when "000001001000"=> s <="100011100001"; -- Argumento 72 Funcion 0.11022221
  when "000001001001"=> s <="100011100100"; -- Argumento 73 Funcion 0.11174671
  when "000001001010"=> s <="100011100111"; -- Argumento 74 Funcion 0.11327095
  when "000001001011"=> s <="100011101011"; -- Argumento 75 Funcion 0.11479493
  when "000001001100"=> s <="100011101110"; -- Argumento 76 Funcion 0.11631863
  when "000001001101"=> s <="100011110001"; -- Argumento 77 Funcion 0.11784206
  when "000001001110"=> s <="100011110100"; -- Argumento 78 Funcion 0.11936521
  when "000001001111"=> s <="100011110111"; -- Argumento 79 Funcion 0.12088809
  when "000001010000"=> s <="100011111010"; -- Argumento 80 Funcion 0.12241068
  when "000001010001"=> s <="100011111101"; -- Argumento 81 Funcion 0.12393298
  when "000001010010"=> s <="100100000000"; -- Argumento 82 Funcion 0.12545498
  when "000001010011"=> s <="100100000100"; -- Argumento 83 Funcion 0.12697670
  when "000001010100"=> s <="100100000111"; -- Argumento 84 Funcion 0.12849811
  when "000001010101"=> s <="100100001010"; -- Argumento 85 Funcion 0.13001922
  when "000001010110"=> s <="100100001101"; -- Argumento 86 Funcion 0.13154003
  when "000001010111"=> s <="100100010000"; -- Argumento 87 Funcion 0.13306053
  when "000001011000"=> s <="100100010011"; -- Argumento 88 Funcion 0.13458071
  when "000001011001"=> s <="100100010110"; -- Argumento 89 Funcion 0.13610058
  when "000001011010"=> s <="100100011001"; -- Argumento 90 Funcion 0.13762012
  when "000001011011"=> s <="100100011100"; -- Argumento 91 Funcion 0.13913934
  when "000001011100"=> s <="100100100000"; -- Argumento 92 Funcion 0.14065824
  when "000001011101"=> s <="100100100011"; -- Argumento 93 Funcion 0.14217680
  when "000001011110"=> s <="100100100110"; -- Argumento 94 Funcion 0.14369503
  when "000001011111"=> s <="100100101001"; -- Argumento 95 Funcion 0.14521292
  when "000001100000"=> s <="100100101100"; -- Argumento 96 Funcion 0.14673047
  when "000001100001"=> s <="100100101111"; -- Argumento 97 Funcion 0.14824768
  when "000001100010"=> s <="100100110010"; -- Argumento 98 Funcion 0.14976453
  when "000001100011"=> s <="100100110101"; -- Argumento 99 Funcion 0.15128104
  when "000001100100"=> s <="100100111000"; -- Argumento 100 Funcion 0.15279719
  when "000001100101"=> s <="100100111100"; -- Argumento 101 Funcion 0.15431297
  when "000001100110"=> s <="100100111111"; -- Argumento 102 Funcion 0.15582840
  when "000001100111"=> s <="100101000010"; -- Argumento 103 Funcion 0.15734346
  when "000001101000"=> s <="100101000101"; -- Argumento 104 Funcion 0.15885814
  when "000001101001"=> s <="100101001000"; -- Argumento 105 Funcion 0.16037246
  when "000001101010"=> s <="100101001011"; -- Argumento 106 Funcion 0.16188639
  when "000001101011"=> s <="100101001110"; -- Argumento 107 Funcion 0.16339995
  when "000001101100"=> s <="100101010001"; -- Argumento 108 Funcion 0.16491312
  when "000001101101"=> s <="100101010100"; -- Argumento 109 Funcion 0.16642590
  when "000001101110"=> s <="100101010111"; -- Argumento 110 Funcion 0.16793829
  when "000001101111"=> s <="100101011011"; -- Argumento 111 Funcion 0.16945029
  when "000001110000"=> s <="100101011110"; -- Argumento 112 Funcion 0.17096189
  when "000001110001"=> s <="100101100001"; -- Argumento 113 Funcion 0.17247308
  when "000001110010"=> s <="100101100100"; -- Argumento 114 Funcion 0.17398387
  when "000001110011"=> s <="100101100111"; -- Argumento 115 Funcion 0.17549425
  when "000001110100"=> s <="100101101010"; -- Argumento 116 Funcion 0.17700422
  when "000001110101"=> s <="100101101101"; -- Argumento 117 Funcion 0.17851377
  when "000001110110"=> s <="100101110000"; -- Argumento 118 Funcion 0.18002290
  when "000001110111"=> s <="100101110011"; -- Argumento 119 Funcion 0.18153161
  when "000001111000"=> s <="100101110110"; -- Argumento 120 Funcion 0.18303989
  when "000001111001"=> s <="100101111001"; -- Argumento 121 Funcion 0.18454774
  when "000001111010"=> s <="100101111101"; -- Argumento 122 Funcion 0.18605515
  when "000001111011"=> s <="100110000000"; -- Argumento 123 Funcion 0.18756213
  when "000001111100"=> s <="100110000011"; -- Argumento 124 Funcion 0.18906866
  when "000001111101"=> s <="100110000110"; -- Argumento 125 Funcion 0.19057475
  when "000001111110"=> s <="100110001001"; -- Argumento 126 Funcion 0.19208040
  when "000001111111"=> s <="100110001100"; -- Argumento 127 Funcion 0.19358559
  when "000010000000"=> s <="100110001111"; -- Argumento 128 Funcion 0.19509032
  when "000010000001"=> s <="100110010010"; -- Argumento 129 Funcion 0.19659460
  when "000010000010"=> s <="100110010101"; -- Argumento 130 Funcion 0.19809841
  when "000010000011"=> s <="100110011000"; -- Argumento 131 Funcion 0.19960176
  when "000010000100"=> s <="100110011011"; -- Argumento 132 Funcion 0.20110463
  when "000010000101"=> s <="100110011110"; -- Argumento 133 Funcion 0.20260704
  when "000010000110"=> s <="100110100010"; -- Argumento 134 Funcion 0.20410897
  when "000010000111"=> s <="100110100101"; -- Argumento 135 Funcion 0.20561041
  when "000010001000"=> s <="100110101000"; -- Argumento 136 Funcion 0.20711138
  when "000010001001"=> s <="100110101011"; -- Argumento 137 Funcion 0.20861185
  when "000010001010"=> s <="100110101110"; -- Argumento 138 Funcion 0.21011184
  when "000010001011"=> s <="100110110001"; -- Argumento 139 Funcion 0.21161133
  when "000010001100"=> s <="100110110100"; -- Argumento 140 Funcion 0.21311032
  when "000010001101"=> s <="100110110111"; -- Argumento 141 Funcion 0.21460881
  when "000010001110"=> s <="100110111010"; -- Argumento 142 Funcion 0.21610680
  when "000010001111"=> s <="100110111101"; -- Argumento 143 Funcion 0.21760427
  when "000010010000"=> s <="100111000000"; -- Argumento 144 Funcion 0.21910124
  when "000010010001"=> s <="100111000011"; -- Argumento 145 Funcion 0.22059769
  when "000010010010"=> s <="100111000110"; -- Argumento 146 Funcion 0.22209362
  when "000010010011"=> s <="100111001001"; -- Argumento 147 Funcion 0.22358903
  when "000010010100"=> s <="100111001100"; -- Argumento 148 Funcion 0.22508391
  when "000010010101"=> s <="100111010000"; -- Argumento 149 Funcion 0.22657826
  when "000010010110"=> s <="100111010011"; -- Argumento 150 Funcion 0.22807208
  when "000010010111"=> s <="100111010110"; -- Argumento 151 Funcion 0.22956537
  when "000010011000"=> s <="100111011001"; -- Argumento 152 Funcion 0.23105811
  when "000010011001"=> s <="100111011100"; -- Argumento 153 Funcion 0.23255031
  when "000010011010"=> s <="100111011111"; -- Argumento 154 Funcion 0.23404196
  when "000010011011"=> s <="100111100010"; -- Argumento 155 Funcion 0.23553306
  when "000010011100"=> s <="100111100101"; -- Argumento 156 Funcion 0.23702361
  when "000010011101"=> s <="100111101000"; -- Argumento 157 Funcion 0.23851359
  when "000010011110"=> s <="100111101011"; -- Argumento 158 Funcion 0.24000302
  when "000010011111"=> s <="100111101110"; -- Argumento 159 Funcion 0.24149189
  when "000010100000"=> s <="100111110001"; -- Argumento 160 Funcion 0.24298018
  when "000010100001"=> s <="100111110100"; -- Argumento 161 Funcion 0.24446790
  when "000010100010"=> s <="100111110111"; -- Argumento 162 Funcion 0.24595505
  when "000010100011"=> s <="100111111010"; -- Argumento 163 Funcion 0.24744162
  when "000010100100"=> s <="100111111101"; -- Argumento 164 Funcion 0.24892761
  when "000010100101"=> s <="101000000000"; -- Argumento 165 Funcion 0.25041301
  when "000010100110"=> s <="101000000011"; -- Argumento 166 Funcion 0.25189782
  when "000010100111"=> s <="101000000110"; -- Argumento 167 Funcion 0.25338204
  when "000010101000"=> s <="101000001001"; -- Argumento 168 Funcion 0.25486566
  when "000010101001"=> s <="101000001101"; -- Argumento 169 Funcion 0.25634868
  when "000010101010"=> s <="101000010000"; -- Argumento 170 Funcion 0.25783110
  when "000010101011"=> s <="101000010011"; -- Argumento 171 Funcion 0.25931292
  when "000010101100"=> s <="101000010110"; -- Argumento 172 Funcion 0.26079412
  when "000010101101"=> s <="101000011001"; -- Argumento 173 Funcion 0.26227471
  when "000010101110"=> s <="101000011100"; -- Argumento 174 Funcion 0.26375468
  when "000010101111"=> s <="101000011111"; -- Argumento 175 Funcion 0.26523403
  when "000010110000"=> s <="101000100010"; -- Argumento 176 Funcion 0.26671276
  when "000010110001"=> s <="101000100101"; -- Argumento 177 Funcion 0.26819086
  when "000010110010"=> s <="101000101000"; -- Argumento 178 Funcion 0.26966833
  when "000010110011"=> s <="101000101011"; -- Argumento 179 Funcion 0.27114516
  when "000010110100"=> s <="101000101110"; -- Argumento 180 Funcion 0.27262136
  when "000010110101"=> s <="101000110001"; -- Argumento 181 Funcion 0.27409691
  when "000010110110"=> s <="101000110100"; -- Argumento 182 Funcion 0.27557182
  when "000010110111"=> s <="101000110111"; -- Argumento 183 Funcion 0.27704608
  when "000010111000"=> s <="101000111010"; -- Argumento 184 Funcion 0.27851969
  when "000010111001"=> s <="101000111101"; -- Argumento 185 Funcion 0.27999264
  when "000010111010"=> s <="101001000000"; -- Argumento 186 Funcion 0.28146494
  when "000010111011"=> s <="101001000011"; -- Argumento 187 Funcion 0.28293657
  when "000010111100"=> s <="101001000110"; -- Argumento 188 Funcion 0.28440754
  when "000010111101"=> s <="101001001001"; -- Argumento 189 Funcion 0.28587783
  when "000010111110"=> s <="101001001100"; -- Argumento 190 Funcion 0.28734746
  when "000010111111"=> s <="101001001111"; -- Argumento 191 Funcion 0.28881641
  when "000011000000"=> s <="101001010010"; -- Argumento 192 Funcion 0.29028468
  when "000011000001"=> s <="101001010101"; -- Argumento 193 Funcion 0.29175226
  when "000011000010"=> s <="101001011000"; -- Argumento 194 Funcion 0.29321916
  when "000011000011"=> s <="101001011011"; -- Argumento 195 Funcion 0.29468537
  when "000011000100"=> s <="101001011110"; -- Argumento 196 Funcion 0.29615089
  when "000011000101"=> s <="101001100001"; -- Argumento 197 Funcion 0.29761571
  when "000011000110"=> s <="101001100100"; -- Argumento 198 Funcion 0.29907983
  when "000011000111"=> s <="101001100111"; -- Argumento 199 Funcion 0.30054324
  when "000011001000"=> s <="101001101010"; -- Argumento 200 Funcion 0.30200595
  when "000011001001"=> s <="101001101101"; -- Argumento 201 Funcion 0.30346795
  when "000011001010"=> s <="101001110000"; -- Argumento 202 Funcion 0.30492923
  when "000011001011"=> s <="101001110011"; -- Argumento 203 Funcion 0.30638980
  when "000011001100"=> s <="101001110110"; -- Argumento 204 Funcion 0.30784964
  when "000011001101"=> s <="101001111001"; -- Argumento 205 Funcion 0.30930876
  when "000011001110"=> s <="101001111100"; -- Argumento 206 Funcion 0.31076715
  when "000011001111"=> s <="101001111111"; -- Argumento 207 Funcion 0.31222481
  when "000011010000"=> s <="101010000010"; -- Argumento 208 Funcion 0.31368174
  when "000011010001"=> s <="101010000101"; -- Argumento 209 Funcion 0.31513793
  when "000011010010"=> s <="101010001000"; -- Argumento 210 Funcion 0.31659338
  when "000011010011"=> s <="101010001011"; -- Argumento 211 Funcion 0.31804808
  when "000011010100"=> s <="101010001110"; -- Argumento 212 Funcion 0.31950203
  when "000011010101"=> s <="101010010001"; -- Argumento 213 Funcion 0.32095523
  when "000011010110"=> s <="101010010100"; -- Argumento 214 Funcion 0.32240768
  when "000011010111"=> s <="101010010111"; -- Argumento 215 Funcion 0.32385937
  when "000011011000"=> s <="101010011010"; -- Argumento 216 Funcion 0.32531029
  when "000011011001"=> s <="101010011101"; -- Argumento 217 Funcion 0.32676045
  when "000011011010"=> s <="101010100000"; -- Argumento 218 Funcion 0.32820984
  when "000011011011"=> s <="101010100011"; -- Argumento 219 Funcion 0.32965846
  when "000011011100"=> s <="101010100110"; -- Argumento 220 Funcion 0.33110631
  when "000011011101"=> s <="101010101001"; -- Argumento 221 Funcion 0.33255337
  when "000011011110"=> s <="101010101100"; -- Argumento 222 Funcion 0.33399965
  when "000011011111"=> s <="101010101110"; -- Argumento 223 Funcion 0.33544515
  when "000011100000"=> s <="101010110001"; -- Argumento 224 Funcion 0.33688985
  when "000011100001"=> s <="101010110100"; -- Argumento 225 Funcion 0.33833377
  when "000011100010"=> s <="101010110111"; -- Argumento 226 Funcion 0.33977688
  when "000011100011"=> s <="101010111010"; -- Argumento 227 Funcion 0.34121920
  when "000011100100"=> s <="101010111101"; -- Argumento 228 Funcion 0.34266072
  when "000011100101"=> s <="101011000000"; -- Argumento 229 Funcion 0.34410143
  when "000011100110"=> s <="101011000011"; -- Argumento 230 Funcion 0.34554132
  when "000011100111"=> s <="101011000110"; -- Argumento 231 Funcion 0.34698041
  when "000011101000"=> s <="101011001001"; -- Argumento 232 Funcion 0.34841868
  when "000011101001"=> s <="101011001100"; -- Argumento 233 Funcion 0.34985613
  when "000011101010"=> s <="101011001111"; -- Argumento 234 Funcion 0.35129276
  when "000011101011"=> s <="101011010010"; -- Argumento 235 Funcion 0.35272856
  when "000011101100"=> s <="101011010101"; -- Argumento 236 Funcion 0.35416353
  when "000011101101"=> s <="101011011000"; -- Argumento 237 Funcion 0.35559766
  when "000011101110"=> s <="101011011011"; -- Argumento 238 Funcion 0.35703096
  when "000011101111"=> s <="101011011110"; -- Argumento 239 Funcion 0.35846342
  when "000011110000"=> s <="101011100001"; -- Argumento 240 Funcion 0.35989504
  when "000011110001"=> s <="101011100011"; -- Argumento 241 Funcion 0.36132581
  when "000011110010"=> s <="101011100110"; -- Argumento 242 Funcion 0.36275572
  when "000011110011"=> s <="101011101001"; -- Argumento 243 Funcion 0.36418479
  when "000011110100"=> s <="101011101100"; -- Argumento 244 Funcion 0.36561300
  when "000011110101"=> s <="101011101111"; -- Argumento 245 Funcion 0.36704035
  when "000011110110"=> s <="101011110010"; -- Argumento 246 Funcion 0.36846683
  when "000011110111"=> s <="101011110101"; -- Argumento 247 Funcion 0.36989245
  when "000011111000"=> s <="101011111000"; -- Argumento 248 Funcion 0.37131719
  when "000011111001"=> s <="101011111011"; -- Argumento 249 Funcion 0.37274107
  when "000011111010"=> s <="101011111110"; -- Argumento 250 Funcion 0.37416406
  when "000011111011"=> s <="101100000001"; -- Argumento 251 Funcion 0.37558618
  when "000011111100"=> s <="101100000100"; -- Argumento 252 Funcion 0.37700741
  when "000011111101"=> s <="101100000111"; -- Argumento 253 Funcion 0.37842775
  when "000011111110"=> s <="101100001001"; -- Argumento 254 Funcion 0.37984721
  when "000011111111"=> s <="101100001100"; -- Argumento 255 Funcion 0.38126577
  when "000100000000"=> s <="101100001111"; -- Argumento 256 Funcion 0.38268343
  when "000100000001"=> s <="101100010010"; -- Argumento 257 Funcion 0.38410020
  when "000100000010"=> s <="101100010101"; -- Argumento 258 Funcion 0.38551605
  when "000100000011"=> s <="101100011000"; -- Argumento 259 Funcion 0.38693101
  when "000100000100"=> s <="101100011011"; -- Argumento 260 Funcion 0.38834505
  when "000100000101"=> s <="101100011110"; -- Argumento 261 Funcion 0.38975817
  when "000100000110"=> s <="101100100001"; -- Argumento 262 Funcion 0.39117038
  when "000100000111"=> s <="101100100100"; -- Argumento 263 Funcion 0.39258167
  when "000100001000"=> s <="101100100110"; -- Argumento 264 Funcion 0.39399204
  when "000100001001"=> s <="101100101001"; -- Argumento 265 Funcion 0.39540148
  when "000100001010"=> s <="101100101100"; -- Argumento 266 Funcion 0.39680999
  when "000100001011"=> s <="101100101111"; -- Argumento 267 Funcion 0.39821756
  when "000100001100"=> s <="101100110010"; -- Argumento 268 Funcion 0.39962420
  when "000100001101"=> s <="101100110101"; -- Argumento 269 Funcion 0.40102990
  when "000100001110"=> s <="101100111000"; -- Argumento 270 Funcion 0.40243465
  when "000100001111"=> s <="101100111011"; -- Argumento 271 Funcion 0.40383846
  when "000100010000"=> s <="101100111101"; -- Argumento 272 Funcion 0.40524131
  when "000100010001"=> s <="101101000000"; -- Argumento 273 Funcion 0.40664322
  when "000100010010"=> s <="101101000011"; -- Argumento 274 Funcion 0.40804416
  when "000100010011"=> s <="101101000110"; -- Argumento 275 Funcion 0.40944415
  when "000100010100"=> s <="101101001001"; -- Argumento 276 Funcion 0.41084317
  when "000100010101"=> s <="101101001100"; -- Argumento 277 Funcion 0.41224123
  when "000100010110"=> s <="101101001111"; -- Argumento 278 Funcion 0.41363831
  when "000100010111"=> s <="101101010001"; -- Argumento 279 Funcion 0.41503442
  when "000100011000"=> s <="101101010100"; -- Argumento 280 Funcion 0.41642956
  when "000100011001"=> s <="101101010111"; -- Argumento 281 Funcion 0.41782372
  when "000100011010"=> s <="101101011010"; -- Argumento 282 Funcion 0.41921689
  when "000100011011"=> s <="101101011101"; -- Argumento 283 Funcion 0.42060907
  when "000100011100"=> s <="101101100000"; -- Argumento 284 Funcion 0.42200027
  when "000100011101"=> s <="101101100011"; -- Argumento 285 Funcion 0.42339047
  when "000100011110"=> s <="101101100101"; -- Argumento 286 Funcion 0.42477968
  when "000100011111"=> s <="101101101000"; -- Argumento 287 Funcion 0.42616789
  when "000100100000"=> s <="101101101011"; -- Argumento 288 Funcion 0.42755509
  when "000100100001"=> s <="101101101110"; -- Argumento 289 Funcion 0.42894129
  when "000100100010"=> s <="101101110001"; -- Argumento 290 Funcion 0.43032648
  when "000100100011"=> s <="101101110100"; -- Argumento 291 Funcion 0.43171066
  when "000100100100"=> s <="101101110110"; -- Argumento 292 Funcion 0.43309382
  when "000100100101"=> s <="101101111001"; -- Argumento 293 Funcion 0.43447596
  when "000100100110"=> s <="101101111100"; -- Argumento 294 Funcion 0.43585708
  when "000100100111"=> s <="101101111111"; -- Argumento 295 Funcion 0.43723717
  when "000100101000"=> s <="101110000010"; -- Argumento 296 Funcion 0.43861624
  when "000100101001"=> s <="101110000101"; -- Argumento 297 Funcion 0.43999427
  when "000100101010"=> s <="101110000111"; -- Argumento 298 Funcion 0.44137127
  when "000100101011"=> s <="101110001010"; -- Argumento 299 Funcion 0.44274723
  when "000100101100"=> s <="101110001101"; -- Argumento 300 Funcion 0.44412214
  when "000100101101"=> s <="101110010000"; -- Argumento 301 Funcion 0.44549602
  when "000100101110"=> s <="101110010011"; -- Argumento 302 Funcion 0.44686884
  when "000100101111"=> s <="101110010101"; -- Argumento 303 Funcion 0.44824061
  when "000100110000"=> s <="101110011000"; -- Argumento 304 Funcion 0.44961133
  when "000100110001"=> s <="101110011011"; -- Argumento 305 Funcion 0.45098099
  when "000100110010"=> s <="101110011110"; -- Argumento 306 Funcion 0.45234959
  when "000100110011"=> s <="101110100001"; -- Argumento 307 Funcion 0.45371712
  when "000100110100"=> s <="101110100100"; -- Argumento 308 Funcion 0.45508359
  when "000100110101"=> s <="101110100110"; -- Argumento 309 Funcion 0.45644898
  when "000100110110"=> s <="101110101001"; -- Argumento 310 Funcion 0.45781330
  when "000100110111"=> s <="101110101100"; -- Argumento 311 Funcion 0.45917655
  when "000100111000"=> s <="101110101111"; -- Argumento 312 Funcion 0.46053871
  when "000100111001"=> s <="101110110001"; -- Argumento 313 Funcion 0.46189979
  when "000100111010"=> s <="101110110100"; -- Argumento 314 Funcion 0.46325978
  when "000100111011"=> s <="101110110111"; -- Argumento 315 Funcion 0.46461869
  when "000100111100"=> s <="101110111010"; -- Argumento 316 Funcion 0.46597650
  when "000100111101"=> s <="101110111101"; -- Argumento 317 Funcion 0.46733321
  when "000100111110"=> s <="101110111111"; -- Argumento 318 Funcion 0.46868882
  when "000100111111"=> s <="101111000010"; -- Argumento 319 Funcion 0.47004333
  when "000101000000"=> s <="101111000101"; -- Argumento 320 Funcion 0.47139674
  when "000101000001"=> s <="101111001000"; -- Argumento 321 Funcion 0.47274903
  when "000101000010"=> s <="101111001010"; -- Argumento 322 Funcion 0.47410021
  when "000101000011"=> s <="101111001101"; -- Argumento 323 Funcion 0.47545028
  when "000101000100"=> s <="101111010000"; -- Argumento 324 Funcion 0.47679923
  when "000101000101"=> s <="101111010011"; -- Argumento 325 Funcion 0.47814706
  when "000101000110"=> s <="101111010110"; -- Argumento 326 Funcion 0.47949376
  when "000101000111"=> s <="101111011000"; -- Argumento 327 Funcion 0.48083933
  when "000101001000"=> s <="101111011011"; -- Argumento 328 Funcion 0.48218377
  when "000101001001"=> s <="101111011110"; -- Argumento 329 Funcion 0.48352708
  when "000101001010"=> s <="101111100001"; -- Argumento 330 Funcion 0.48486925
  when "000101001011"=> s <="101111100011"; -- Argumento 331 Funcion 0.48621028
  when "000101001100"=> s <="101111100110"; -- Argumento 332 Funcion 0.48755016
  when "000101001101"=> s <="101111101001"; -- Argumento 333 Funcion 0.48888890
  when "000101001110"=> s <="101111101011"; -- Argumento 334 Funcion 0.49022648
  when "000101001111"=> s <="101111101110"; -- Argumento 335 Funcion 0.49156292
  when "000101010000"=> s <="101111110001"; -- Argumento 336 Funcion 0.49289819
  when "000101010001"=> s <="101111110100"; -- Argumento 337 Funcion 0.49423231
  when "000101010010"=> s <="101111110110"; -- Argumento 338 Funcion 0.49556526
  when "000101010011"=> s <="101111111001"; -- Argumento 339 Funcion 0.49689705
  when "000101010100"=> s <="101111111100"; -- Argumento 340 Funcion 0.49822767
  when "000101010101"=> s <="101111111111"; -- Argumento 341 Funcion 0.49955711
  when "000101010110"=> s <="110000000001"; -- Argumento 342 Funcion 0.50088538
  when "000101010111"=> s <="110000000100"; -- Argumento 343 Funcion 0.50221247
  when "000101011000"=> s <="110000000111"; -- Argumento 344 Funcion 0.50353838
  when "000101011001"=> s <="110000001001"; -- Argumento 345 Funcion 0.50486311
  when "000101011010"=> s <="110000001100"; -- Argumento 346 Funcion 0.50618665
  when "000101011011"=> s <="110000001111"; -- Argumento 347 Funcion 0.50750899
  when "000101011100"=> s <="110000010010"; -- Argumento 348 Funcion 0.50883014
  when "000101011101"=> s <="110000010100"; -- Argumento 349 Funcion 0.51015010
  when "000101011110"=> s <="110000010111"; -- Argumento 350 Funcion 0.51146885
  when "000101011111"=> s <="110000011010"; -- Argumento 351 Funcion 0.51278640
  when "000101100000"=> s <="110000011100"; -- Argumento 352 Funcion 0.51410274
  when "000101100001"=> s <="110000011111"; -- Argumento 353 Funcion 0.51541788
  when "000101100010"=> s <="110000100010"; -- Argumento 354 Funcion 0.51673180
  when "000101100011"=> s <="110000100100"; -- Argumento 355 Funcion 0.51804450
  when "000101100100"=> s <="110000100111"; -- Argumento 356 Funcion 0.51935599
  when "000101100101"=> s <="110000101010"; -- Argumento 357 Funcion 0.52066625
  when "000101100110"=> s <="110000101101"; -- Argumento 358 Funcion 0.52197529
  when "000101100111"=> s <="110000101111"; -- Argumento 359 Funcion 0.52328310
  when "000101101000"=> s <="110000110010"; -- Argumento 360 Funcion 0.52458968
  when "000101101001"=> s <="110000110101"; -- Argumento 361 Funcion 0.52589503
  when "000101101010"=> s <="110000110111"; -- Argumento 362 Funcion 0.52719913
  when "000101101011"=> s <="110000111010"; -- Argumento 363 Funcion 0.52850200
  when "000101101100"=> s <="110000111101"; -- Argumento 364 Funcion 0.52980362
  when "000101101101"=> s <="110000111111"; -- Argumento 365 Funcion 0.53110400
  when "000101101110"=> s <="110001000010"; -- Argumento 366 Funcion 0.53240313
  when "000101101111"=> s <="110001000101"; -- Argumento 367 Funcion 0.53370100
  when "000101110000"=> s <="110001000111"; -- Argumento 368 Funcion 0.53499762
  when "000101110001"=> s <="110001001010"; -- Argumento 369 Funcion 0.53629298
  when "000101110010"=> s <="110001001100"; -- Argumento 370 Funcion 0.53758708
  when "000101110011"=> s <="110001001111"; -- Argumento 371 Funcion 0.53887991
  when "000101110100"=> s <="110001010010"; -- Argumento 372 Funcion 0.54017147
  when "000101110101"=> s <="110001010100"; -- Argumento 373 Funcion 0.54146177
  when "000101110110"=> s <="110001010111"; -- Argumento 374 Funcion 0.54275078
  when "000101110111"=> s <="110001011010"; -- Argumento 375 Funcion 0.54403853
  when "000101111000"=> s <="110001011100"; -- Argumento 376 Funcion 0.54532499
  when "000101111001"=> s <="110001011111"; -- Argumento 377 Funcion 0.54661017
  when "000101111010"=> s <="110001100010"; -- Argumento 378 Funcion 0.54789406
  when "000101111011"=> s <="110001100100"; -- Argumento 379 Funcion 0.54917666
  when "000101111100"=> s <="110001100111"; -- Argumento 380 Funcion 0.55045797
  when "000101111101"=> s <="110001101001"; -- Argumento 381 Funcion 0.55173799
  when "000101111110"=> s <="110001101100"; -- Argumento 382 Funcion 0.55301671
  when "000101111111"=> s <="110001101111"; -- Argumento 383 Funcion 0.55429412
  when "000110000000"=> s <="110001110001"; -- Argumento 384 Funcion 0.55557023
  when "000110000001"=> s <="110001110100"; -- Argumento 385 Funcion 0.55684504
  when "000110000010"=> s <="110001110111"; -- Argumento 386 Funcion 0.55811853
  when "000110000011"=> s <="110001111001"; -- Argumento 387 Funcion 0.55939071
  when "000110000100"=> s <="110001111100"; -- Argumento 388 Funcion 0.56066158
  when "000110000101"=> s <="110001111110"; -- Argumento 389 Funcion 0.56193112
  when "000110000110"=> s <="110010000001"; -- Argumento 390 Funcion 0.56319934
  when "000110000111"=> s <="110010000100"; -- Argumento 391 Funcion 0.56446624
  when "000110001000"=> s <="110010000110"; -- Argumento 392 Funcion 0.56573181
  when "000110001001"=> s <="110010001001"; -- Argumento 393 Funcion 0.56699605
  when "000110001010"=> s <="110010001011"; -- Argumento 394 Funcion 0.56825895
  when "000110001011"=> s <="110010001110"; -- Argumento 395 Funcion 0.56952052
  when "000110001100"=> s <="110010010000"; -- Argumento 396 Funcion 0.57078075
  when "000110001101"=> s <="110010010011"; -- Argumento 397 Funcion 0.57203963
  when "000110001110"=> s <="110010010110"; -- Argumento 398 Funcion 0.57329717
  when "000110001111"=> s <="110010011000"; -- Argumento 399 Funcion 0.57455336
  when "000110010000"=> s <="110010011011"; -- Argumento 400 Funcion 0.57580819
  when "000110010001"=> s <="110010011101"; -- Argumento 401 Funcion 0.57706167
  when "000110010010"=> s <="110010100000"; -- Argumento 402 Funcion 0.57831380
  when "000110010011"=> s <="110010100010"; -- Argumento 403 Funcion 0.57956456
  when "000110010100"=> s <="110010100101"; -- Argumento 404 Funcion 0.58081396
  when "000110010101"=> s <="110010101000"; -- Argumento 405 Funcion 0.58206199
  when "000110010110"=> s <="110010101010"; -- Argumento 406 Funcion 0.58330865
  when "000110010111"=> s <="110010101101"; -- Argumento 407 Funcion 0.58455394
  when "000110011000"=> s <="110010101111"; -- Argumento 408 Funcion 0.58579786
  when "000110011001"=> s <="110010110010"; -- Argumento 409 Funcion 0.58704039
  when "000110011010"=> s <="110010110100"; -- Argumento 410 Funcion 0.58828155
  when "000110011011"=> s <="110010110111"; -- Argumento 411 Funcion 0.58952132
  when "000110011100"=> s <="110010111001"; -- Argumento 412 Funcion 0.59075970
  when "000110011101"=> s <="110010111100"; -- Argumento 413 Funcion 0.59199669
  when "000110011110"=> s <="110010111110"; -- Argumento 414 Funcion 0.59323230
  when "000110011111"=> s <="110011000001"; -- Argumento 415 Funcion 0.59446650
  when "000110100000"=> s <="110011000011"; -- Argumento 416 Funcion 0.59569930
  when "000110100001"=> s <="110011000110"; -- Argumento 417 Funcion 0.59693071
  when "000110100010"=> s <="110011001001"; -- Argumento 418 Funcion 0.59816071
  when "000110100011"=> s <="110011001011"; -- Argumento 419 Funcion 0.59938930
  when "000110100100"=> s <="110011001110"; -- Argumento 420 Funcion 0.60061648
  when "000110100101"=> s <="110011010000"; -- Argumento 421 Funcion 0.60184225
  when "000110100110"=> s <="110011010011"; -- Argumento 422 Funcion 0.60306660
  when "000110100111"=> s <="110011010101"; -- Argumento 423 Funcion 0.60428953
  when "000110101000"=> s <="110011011000"; -- Argumento 424 Funcion 0.60551104
  when "000110101001"=> s <="110011011010"; -- Argumento 425 Funcion 0.60673113
  when "000110101010"=> s <="110011011101"; -- Argumento 426 Funcion 0.60794978
  when "000110101011"=> s <="110011011111"; -- Argumento 427 Funcion 0.60916701
  when "000110101100"=> s <="110011100010"; -- Argumento 428 Funcion 0.61038281
  when "000110101101"=> s <="110011100100"; -- Argumento 429 Funcion 0.61159716
  when "000110101110"=> s <="110011100111"; -- Argumento 430 Funcion 0.61281008
  when "000110101111"=> s <="110011101001"; -- Argumento 431 Funcion 0.61402156
  when "000110110000"=> s <="110011101011"; -- Argumento 432 Funcion 0.61523159
  when "000110110001"=> s <="110011101110"; -- Argumento 433 Funcion 0.61644017
  when "000110110010"=> s <="110011110000"; -- Argumento 434 Funcion 0.61764731
  when "000110110011"=> s <="110011110011"; -- Argumento 435 Funcion 0.61885299
  when "000110110100"=> s <="110011110101"; -- Argumento 436 Funcion 0.62005721
  when "000110110101"=> s <="110011111000"; -- Argumento 437 Funcion 0.62125998
  when "000110110110"=> s <="110011111010"; -- Argumento 438 Funcion 0.62246128
  when "000110110111"=> s <="110011111101"; -- Argumento 439 Funcion 0.62366112
  when "000110111000"=> s <="110011111111"; -- Argumento 440 Funcion 0.62485949
  when "000110111001"=> s <="110100000010"; -- Argumento 441 Funcion 0.62605639
  when "000110111010"=> s <="110100000100"; -- Argumento 442 Funcion 0.62725182
  when "000110111011"=> s <="110100000111"; -- Argumento 443 Funcion 0.62844577
  when "000110111100"=> s <="110100001001"; -- Argumento 444 Funcion 0.62963824
  when "000110111101"=> s <="110100001011"; -- Argumento 445 Funcion 0.63082923
  when "000110111110"=> s <="110100001110"; -- Argumento 446 Funcion 0.63201874
  when "000110111111"=> s <="110100010000"; -- Argumento 447 Funcion 0.63320676
  when "000111000000"=> s <="110100010011"; -- Argumento 448 Funcion 0.63439328
  when "000111000001"=> s <="110100010101"; -- Argumento 449 Funcion 0.63557832
  when "000111000010"=> s <="110100011000"; -- Argumento 450 Funcion 0.63676186
  when "000111000011"=> s <="110100011010"; -- Argumento 451 Funcion 0.63794390
  when "000111000100"=> s <="110100011100"; -- Argumento 452 Funcion 0.63912444
  when "000111000101"=> s <="110100011111"; -- Argumento 453 Funcion 0.64030348
  when "000111000110"=> s <="110100100001"; -- Argumento 454 Funcion 0.64148101
  when "000111000111"=> s <="110100100100"; -- Argumento 455 Funcion 0.64265703
  when "000111001000"=> s <="110100100110"; -- Argumento 456 Funcion 0.64383154
  when "000111001001"=> s <="110100101000"; -- Argumento 457 Funcion 0.64500454
  when "000111001010"=> s <="110100101011"; -- Argumento 458 Funcion 0.64617601
  when "000111001011"=> s <="110100101101"; -- Argumento 459 Funcion 0.64734597
  when "000111001100"=> s <="110100110000"; -- Argumento 460 Funcion 0.64851440
  when "000111001101"=> s <="110100110010"; -- Argumento 461 Funcion 0.64968131
  when "000111001110"=> s <="110100110100"; -- Argumento 462 Funcion 0.65084668
  when "000111001111"=> s <="110100110111"; -- Argumento 463 Funcion 0.65201053
  when "000111010000"=> s <="110100111001"; -- Argumento 464 Funcion 0.65317284
  when "000111010001"=> s <="110100111100"; -- Argumento 465 Funcion 0.65433362
  when "000111010010"=> s <="110100111110"; -- Argumento 466 Funcion 0.65549285
  when "000111010011"=> s <="110101000000"; -- Argumento 467 Funcion 0.65665055
  when "000111010100"=> s <="110101000011"; -- Argumento 468 Funcion 0.65780669
  when "000111010101"=> s <="110101000101"; -- Argumento 469 Funcion 0.65896129
  when "000111010110"=> s <="110101000111"; -- Argumento 470 Funcion 0.66011434
  when "000111010111"=> s <="110101001010"; -- Argumento 471 Funcion 0.66126584
  when "000111011000"=> s <="110101001100"; -- Argumento 472 Funcion 0.66241578
  when "000111011001"=> s <="110101001110"; -- Argumento 473 Funcion 0.66356416
  when "000111011010"=> s <="110101010001"; -- Argumento 474 Funcion 0.66471098
  when "000111011011"=> s <="110101010011"; -- Argumento 475 Funcion 0.66585623
  when "000111011100"=> s <="110101010110"; -- Argumento 476 Funcion 0.66699992
  when "000111011101"=> s <="110101011000"; -- Argumento 477 Funcion 0.66814204
  when "000111011110"=> s <="110101011010"; -- Argumento 478 Funcion 0.66928259
  when "000111011111"=> s <="110101011101"; -- Argumento 479 Funcion 0.67042156
  when "000111100000"=> s <="110101011111"; -- Argumento 480 Funcion 0.67155895
  when "000111100001"=> s <="110101100001"; -- Argumento 481 Funcion 0.67269477
  when "000111100010"=> s <="110101100100"; -- Argumento 482 Funcion 0.67382900
  when "000111100011"=> s <="110101100110"; -- Argumento 483 Funcion 0.67496165
  when "000111100100"=> s <="110101101000"; -- Argumento 484 Funcion 0.67609270
  when "000111100101"=> s <="110101101010"; -- Argumento 485 Funcion 0.67722217
  when "000111100110"=> s <="110101101101"; -- Argumento 486 Funcion 0.67835004
  when "000111100111"=> s <="110101101111"; -- Argumento 487 Funcion 0.67947632
  when "000111101000"=> s <="110101110001"; -- Argumento 488 Funcion 0.68060100
  when "000111101001"=> s <="110101110100"; -- Argumento 489 Funcion 0.68172407
  when "000111101010"=> s <="110101110110"; -- Argumento 490 Funcion 0.68284555
  when "000111101011"=> s <="110101111000"; -- Argumento 491 Funcion 0.68396541
  when "000111101100"=> s <="110101111011"; -- Argumento 492 Funcion 0.68508367
  when "000111101101"=> s <="110101111101"; -- Argumento 493 Funcion 0.68620031
  when "000111101110"=> s <="110101111111"; -- Argumento 494 Funcion 0.68731534
  when "000111101111"=> s <="110110000001"; -- Argumento 495 Funcion 0.68842875
  when "000111110000"=> s <="110110000100"; -- Argumento 496 Funcion 0.68954054
  when "000111110001"=> s <="110110000110"; -- Argumento 497 Funcion 0.69065071
  when "000111110010"=> s <="110110001000"; -- Argumento 498 Funcion 0.69175926
  when "000111110011"=> s <="110110001010"; -- Argumento 499 Funcion 0.69286617
  when "000111110100"=> s <="110110001101"; -- Argumento 500 Funcion 0.69397146
  when "000111110101"=> s <="110110001111"; -- Argumento 501 Funcion 0.69507511
  when "000111110110"=> s <="110110010001"; -- Argumento 502 Funcion 0.69617713
  when "000111110111"=> s <="110110010100"; -- Argumento 503 Funcion 0.69727751
  when "000111111000"=> s <="110110010110"; -- Argumento 504 Funcion 0.69837625
  when "000111111001"=> s <="110110011000"; -- Argumento 505 Funcion 0.69947334
  when "000111111010"=> s <="110110011010"; -- Argumento 506 Funcion 0.70056879
  when "000111111011"=> s <="110110011101"; -- Argumento 507 Funcion 0.70166259
  when "000111111100"=> s <="110110011111"; -- Argumento 508 Funcion 0.70275474
  when "000111111101"=> s <="110110100001"; -- Argumento 509 Funcion 0.70384524
  when "000111111110"=> s <="110110100011"; -- Argumento 510 Funcion 0.70493408
  when "000111111111"=> s <="110110100101"; -- Argumento 511 Funcion 0.70602126
  when "001000000000"=> s <="110110101000"; -- Argumento 512 Funcion 0.70710678
  when "001000000001"=> s <="110110101010"; -- Argumento 513 Funcion 0.70819064
  when "001000000010"=> s <="110110101100"; -- Argumento 514 Funcion 0.70927283
  when "001000000011"=> s <="110110101110"; -- Argumento 515 Funcion 0.71035335
  when "001000000100"=> s <="110110110001"; -- Argumento 516 Funcion 0.71143220
  when "001000000101"=> s <="110110110011"; -- Argumento 517 Funcion 0.71250937
  when "001000000110"=> s <="110110110101"; -- Argumento 518 Funcion 0.71358487
  when "001000000111"=> s <="110110110111"; -- Argumento 519 Funcion 0.71465869
  when "001000001000"=> s <="110110111001"; -- Argumento 520 Funcion 0.71573083
  when "001000001001"=> s <="110110111100"; -- Argumento 521 Funcion 0.71680128
  when "001000001010"=> s <="110110111110"; -- Argumento 522 Funcion 0.71787005
  when "001000001011"=> s <="110111000000"; -- Argumento 523 Funcion 0.71893712
  when "001000001100"=> s <="110111000010"; -- Argumento 524 Funcion 0.72000251
  when "001000001101"=> s <="110111000100"; -- Argumento 525 Funcion 0.72106620
  when "001000001110"=> s <="110111000110"; -- Argumento 526 Funcion 0.72212819
  when "001000001111"=> s <="110111001001"; -- Argumento 527 Funcion 0.72318849
  when "001000010000"=> s <="110111001011"; -- Argumento 528 Funcion 0.72424708
  when "001000010001"=> s <="110111001101"; -- Argumento 529 Funcion 0.72530397
  when "001000010010"=> s <="110111001111"; -- Argumento 530 Funcion 0.72635916
  when "001000010011"=> s <="110111010001"; -- Argumento 531 Funcion 0.72741263
  when "001000010100"=> s <="110111010011"; -- Argumento 532 Funcion 0.72846439
  when "001000010101"=> s <="110111010110"; -- Argumento 533 Funcion 0.72951444
  when "001000010110"=> s <="110111011000"; -- Argumento 534 Funcion 0.73056277
  when "001000010111"=> s <="110111011010"; -- Argumento 535 Funcion 0.73160938
  when "001000011000"=> s <="110111011100"; -- Argumento 536 Funcion 0.73265427
  when "001000011001"=> s <="110111011110"; -- Argumento 537 Funcion 0.73369744
  when "001000011010"=> s <="110111100000"; -- Argumento 538 Funcion 0.73473888
  when "001000011011"=> s <="110111100010"; -- Argumento 539 Funcion 0.73577859
  when "001000011100"=> s <="110111100101"; -- Argumento 540 Funcion 0.73681657
  when "001000011101"=> s <="110111100111"; -- Argumento 541 Funcion 0.73785281
  when "001000011110"=> s <="110111101001"; -- Argumento 542 Funcion 0.73888732
  when "001000011111"=> s <="110111101011"; -- Argumento 543 Funcion 0.73992010
  when "001000100000"=> s <="110111101101"; -- Argumento 544 Funcion 0.74095113
  when "001000100001"=> s <="110111101111"; -- Argumento 545 Funcion 0.74198041
  when "001000100010"=> s <="110111110001"; -- Argumento 546 Funcion 0.74300795
  when "001000100011"=> s <="110111110011"; -- Argumento 547 Funcion 0.74403374
  when "001000100100"=> s <="110111110101"; -- Argumento 548 Funcion 0.74505779
  when "001000100101"=> s <="110111110111"; -- Argumento 549 Funcion 0.74608007
  when "001000100110"=> s <="110111111010"; -- Argumento 550 Funcion 0.74710061
  when "001000100111"=> s <="110111111100"; -- Argumento 551 Funcion 0.74811938
  when "001000101000"=> s <="110111111110"; -- Argumento 552 Funcion 0.74913639
  when "001000101001"=> s <="111000000000"; -- Argumento 553 Funcion 0.75015165
  when "001000101010"=> s <="111000000010"; -- Argumento 554 Funcion 0.75116513
  when "001000101011"=> s <="111000000100"; -- Argumento 555 Funcion 0.75217685
  when "001000101100"=> s <="111000000110"; -- Argumento 556 Funcion 0.75318680
  when "001000101101"=> s <="111000001000"; -- Argumento 557 Funcion 0.75419498
  when "001000101110"=> s <="111000001010"; -- Argumento 558 Funcion 0.75520138
  when "001000101111"=> s <="111000001100"; -- Argumento 559 Funcion 0.75620600
  when "001000110000"=> s <="111000001110"; -- Argumento 560 Funcion 0.75720885
  when "001000110001"=> s <="111000010000"; -- Argumento 561 Funcion 0.75820991
  when "001000110010"=> s <="111000010010"; -- Argumento 562 Funcion 0.75920919
  when "001000110011"=> s <="111000010100"; -- Argumento 563 Funcion 0.76020668
  when "001000110100"=> s <="111000010110"; -- Argumento 564 Funcion 0.76120239
  when "001000110101"=> s <="111000011000"; -- Argumento 565 Funcion 0.76219630
  when "001000110110"=> s <="111000011011"; -- Argumento 566 Funcion 0.76318842
  when "001000110111"=> s <="111000011101"; -- Argumento 567 Funcion 0.76417874
  when "001000111000"=> s <="111000011111"; -- Argumento 568 Funcion 0.76516727
  when "001000111001"=> s <="111000100001"; -- Argumento 569 Funcion 0.76615399
  when "001000111010"=> s <="111000100011"; -- Argumento 570 Funcion 0.76713891
  when "001000111011"=> s <="111000100101"; -- Argumento 571 Funcion 0.76812203
  when "001000111100"=> s <="111000100111"; -- Argumento 572 Funcion 0.76910334
  when "001000111101"=> s <="111000101001"; -- Argumento 573 Funcion 0.77008284
  when "001000111110"=> s <="111000101011"; -- Argumento 574 Funcion 0.77106052
  when "001000111111"=> s <="111000101101"; -- Argumento 575 Funcion 0.77203640
  when "001001000000"=> s <="111000101111"; -- Argumento 576 Funcion 0.77301045
  when "001001000001"=> s <="111000110001"; -- Argumento 577 Funcion 0.77398269
  when "001001000010"=> s <="111000110011"; -- Argumento 578 Funcion 0.77495311
  when "001001000011"=> s <="111000110101"; -- Argumento 579 Funcion 0.77592170
  when "001001000100"=> s <="111000110111"; -- Argumento 580 Funcion 0.77688847
  when "001001000101"=> s <="111000111001"; -- Argumento 581 Funcion 0.77785340
  when "001001000110"=> s <="111000111011"; -- Argumento 582 Funcion 0.77881651
  when "001001000111"=> s <="111000111100"; -- Argumento 583 Funcion 0.77977779
  when "001001001000"=> s <="111000111110"; -- Argumento 584 Funcion 0.78073723
  when "001001001001"=> s <="111001000000"; -- Argumento 585 Funcion 0.78169483
  when "001001001010"=> s <="111001000010"; -- Argumento 586 Funcion 0.78265060
  when "001001001011"=> s <="111001000100"; -- Argumento 587 Funcion 0.78360452
  when "001001001100"=> s <="111001000110"; -- Argumento 588 Funcion 0.78455660
  when "001001001101"=> s <="111001001000"; -- Argumento 589 Funcion 0.78550683
  when "001001001110"=> s <="111001001010"; -- Argumento 590 Funcion 0.78645521
  when "001001001111"=> s <="111001001100"; -- Argumento 591 Funcion 0.78740175
  when "001001010000"=> s <="111001001110"; -- Argumento 592 Funcion 0.78834643
  when "001001010001"=> s <="111001010000"; -- Argumento 593 Funcion 0.78928925
  when "001001010010"=> s <="111001010010"; -- Argumento 594 Funcion 0.79023022
  when "001001010011"=> s <="111001010100"; -- Argumento 595 Funcion 0.79116933
  when "001001010100"=> s <="111001010110"; -- Argumento 596 Funcion 0.79210658
  when "001001010101"=> s <="111001011000"; -- Argumento 597 Funcion 0.79304196
  when "001001010110"=> s <="111001011010"; -- Argumento 598 Funcion 0.79397548
  when "001001010111"=> s <="111001011011"; -- Argumento 599 Funcion 0.79490713
  when "001001011000"=> s <="111001011101"; -- Argumento 600 Funcion 0.79583690
  when "001001011001"=> s <="111001011111"; -- Argumento 601 Funcion 0.79676481
  when "001001011010"=> s <="111001100001"; -- Argumento 602 Funcion 0.79769084
  when "001001011011"=> s <="111001100011"; -- Argumento 603 Funcion 0.79861499
  when "001001011100"=> s <="111001100101"; -- Argumento 604 Funcion 0.79953727
  when "001001011101"=> s <="111001100111"; -- Argumento 605 Funcion 0.80045766
  when "001001011110"=> s <="111001101001"; -- Argumento 606 Funcion 0.80137617
  when "001001011111"=> s <="111001101011"; -- Argumento 607 Funcion 0.80229280
  when "001001100000"=> s <="111001101100"; -- Argumento 608 Funcion 0.80320753
  when "001001100001"=> s <="111001101110"; -- Argumento 609 Funcion 0.80412038
  when "001001100010"=> s <="111001110000"; -- Argumento 610 Funcion 0.80503133
  when "001001100011"=> s <="111001110010"; -- Argumento 611 Funcion 0.80594039
  when "001001100100"=> s <="111001110100"; -- Argumento 612 Funcion 0.80684755
  when "001001100101"=> s <="111001110110"; -- Argumento 613 Funcion 0.80775282
  when "001001100110"=> s <="111001111000"; -- Argumento 614 Funcion 0.80865618
  when "001001100111"=> s <="111001111001"; -- Argumento 615 Funcion 0.80955764
  when "001001101000"=> s <="111001111011"; -- Argumento 616 Funcion 0.81045720
  when "001001101001"=> s <="111001111101"; -- Argumento 617 Funcion 0.81135485
  when "001001101010"=> s <="111001111111"; -- Argumento 618 Funcion 0.81225059
  when "001001101011"=> s <="111010000001"; -- Argumento 619 Funcion 0.81314441
  when "001001101100"=> s <="111010000011"; -- Argumento 620 Funcion 0.81403633
  when "001001101101"=> s <="111010000100"; -- Argumento 621 Funcion 0.81492633
  when "001001101110"=> s <="111010000110"; -- Argumento 622 Funcion 0.81581441
  when "001001101111"=> s <="111010001000"; -- Argumento 623 Funcion 0.81670057
  when "001001110000"=> s <="111010001010"; -- Argumento 624 Funcion 0.81758481
  when "001001110001"=> s <="111010001100"; -- Argumento 625 Funcion 0.81846713
  when "001001110010"=> s <="111010001110"; -- Argumento 626 Funcion 0.81934752
  when "001001110011"=> s <="111010001111"; -- Argumento 627 Funcion 0.82022598
  when "001001110100"=> s <="111010010001"; -- Argumento 628 Funcion 0.82110251
  when "001001110101"=> s <="111010010011"; -- Argumento 629 Funcion 0.82197712
  when "001001110110"=> s <="111010010101"; -- Argumento 630 Funcion 0.82284978
  when "001001110111"=> s <="111010010110"; -- Argumento 631 Funcion 0.82372051
  when "001001111000"=> s <="111010011000"; -- Argumento 632 Funcion 0.82458930
  when "001001111001"=> s <="111010011010"; -- Argumento 633 Funcion 0.82545615
  when "001001111010"=> s <="111010011100"; -- Argumento 634 Funcion 0.82632106
  when "001001111011"=> s <="111010011110"; -- Argumento 635 Funcion 0.82718403
  when "001001111100"=> s <="111010011111"; -- Argumento 636 Funcion 0.82804505
  when "001001111101"=> s <="111010100001"; -- Argumento 637 Funcion 0.82890411
  when "001001111110"=> s <="111010100011"; -- Argumento 638 Funcion 0.82976123
  when "001001111111"=> s <="111010100101"; -- Argumento 639 Funcion 0.83061640
  when "001010000000"=> s <="111010100110"; -- Argumento 640 Funcion 0.83146961
  when "001010000001"=> s <="111010101000"; -- Argumento 641 Funcion 0.83232087
  when "001010000010"=> s <="111010101010"; -- Argumento 642 Funcion 0.83317016
  when "001010000011"=> s <="111010101100"; -- Argumento 643 Funcion 0.83401750
  when "001010000100"=> s <="111010101101"; -- Argumento 644 Funcion 0.83486287
  when "001010000101"=> s <="111010101111"; -- Argumento 645 Funcion 0.83570628
  when "001010000110"=> s <="111010110001"; -- Argumento 646 Funcion 0.83654773
  when "001010000111"=> s <="111010110010"; -- Argumento 647 Funcion 0.83738720
  when "001010001000"=> s <="111010110100"; -- Argumento 648 Funcion 0.83822471
  when "001010001001"=> s <="111010110110"; -- Argumento 649 Funcion 0.83906024
  when "001010001010"=> s <="111010111000"; -- Argumento 650 Funcion 0.83989379
  when "001010001011"=> s <="111010111001"; -- Argumento 651 Funcion 0.84072537
  when "001010001100"=> s <="111010111011"; -- Argumento 652 Funcion 0.84155498
  when "001010001101"=> s <="111010111101"; -- Argumento 653 Funcion 0.84238260
  when "001010001110"=> s <="111010111110"; -- Argumento 654 Funcion 0.84320824
  when "001010001111"=> s <="111011000000"; -- Argumento 655 Funcion 0.84403190
  when "001010010000"=> s <="111011000010"; -- Argumento 656 Funcion 0.84485357
  when "001010010001"=> s <="111011000011"; -- Argumento 657 Funcion 0.84567325
  when "001010010010"=> s <="111011000101"; -- Argumento 658 Funcion 0.84649094
  when "001010010011"=> s <="111011000111"; -- Argumento 659 Funcion 0.84730664
  when "001010010100"=> s <="111011001000"; -- Argumento 660 Funcion 0.84812034
  when "001010010101"=> s <="111011001010"; -- Argumento 661 Funcion 0.84893206
  when "001010010110"=> s <="111011001100"; -- Argumento 662 Funcion 0.84974177
  when "001010010111"=> s <="111011001101"; -- Argumento 663 Funcion 0.85054948
  when "001010011000"=> s <="111011001111"; -- Argumento 664 Funcion 0.85135519
  when "001010011001"=> s <="111011010001"; -- Argumento 665 Funcion 0.85215890
  when "001010011010"=> s <="111011010010"; -- Argumento 666 Funcion 0.85296060
  when "001010011011"=> s <="111011010100"; -- Argumento 667 Funcion 0.85376030
  when "001010011100"=> s <="111011010110"; -- Argumento 668 Funcion 0.85455799
  when "001010011101"=> s <="111011010111"; -- Argumento 669 Funcion 0.85535366
  when "001010011110"=> s <="111011011001"; -- Argumento 670 Funcion 0.85614733
  when "001010011111"=> s <="111011011011"; -- Argumento 671 Funcion 0.85693898
  when "001010100000"=> s <="111011011100"; -- Argumento 672 Funcion 0.85772861
  when "001010100001"=> s <="111011011110"; -- Argumento 673 Funcion 0.85851622
  when "001010100010"=> s <="111011011111"; -- Argumento 674 Funcion 0.85930182
  when "001010100011"=> s <="111011100001"; -- Argumento 675 Funcion 0.86008539
  when "001010100100"=> s <="111011100011"; -- Argumento 676 Funcion 0.86086694
  when "001010100101"=> s <="111011100100"; -- Argumento 677 Funcion 0.86164646
  when "001010100110"=> s <="111011100110"; -- Argumento 678 Funcion 0.86242396
  when "001010100111"=> s <="111011100111"; -- Argumento 679 Funcion 0.86319942
  when "001010101000"=> s <="111011101001"; -- Argumento 680 Funcion 0.86397286
  when "001010101001"=> s <="111011101010"; -- Argumento 681 Funcion 0.86474426
  when "001010101010"=> s <="111011101100"; -- Argumento 682 Funcion 0.86551362
  when "001010101011"=> s <="111011101110"; -- Argumento 683 Funcion 0.86628095
  when "001010101100"=> s <="111011101111"; -- Argumento 684 Funcion 0.86704625
  when "001010101101"=> s <="111011110001"; -- Argumento 685 Funcion 0.86780950
  when "001010101110"=> s <="111011110010"; -- Argumento 686 Funcion 0.86857071
  when "001010101111"=> s <="111011110100"; -- Argumento 687 Funcion 0.86932987
  when "001010110000"=> s <="111011110101"; -- Argumento 688 Funcion 0.87008699
  when "001010110001"=> s <="111011110111"; -- Argumento 689 Funcion 0.87084206
  when "001010110010"=> s <="111011111001"; -- Argumento 690 Funcion 0.87159509
  when "001010110011"=> s <="111011111010"; -- Argumento 691 Funcion 0.87234606
  when "001010110100"=> s <="111011111100"; -- Argumento 692 Funcion 0.87309498
  when "001010110101"=> s <="111011111101"; -- Argumento 693 Funcion 0.87384184
  when "001010110110"=> s <="111011111111"; -- Argumento 694 Funcion 0.87458665
  when "001010110111"=> s <="111100000000"; -- Argumento 695 Funcion 0.87532940
  when "001010111000"=> s <="111100000010"; -- Argumento 696 Funcion 0.87607009
  when "001010111001"=> s <="111100000011"; -- Argumento 697 Funcion 0.87680872
  when "001010111010"=> s <="111100000101"; -- Argumento 698 Funcion 0.87754529
  when "001010111011"=> s <="111100000110"; -- Argumento 699 Funcion 0.87827979
  when "001010111100"=> s <="111100001000"; -- Argumento 700 Funcion 0.87901223
  when "001010111101"=> s <="111100001001"; -- Argumento 701 Funcion 0.87974259
  when "001010111110"=> s <="111100001011"; -- Argumento 702 Funcion 0.88047089
  when "001010111111"=> s <="111100001100"; -- Argumento 703 Funcion 0.88119711
  when "001011000000"=> s <="111100001110"; -- Argumento 704 Funcion 0.88192126
  when "001011000001"=> s <="111100001111"; -- Argumento 705 Funcion 0.88264334
  when "001011000010"=> s <="111100010001"; -- Argumento 706 Funcion 0.88336334
  when "001011000011"=> s <="111100010010"; -- Argumento 707 Funcion 0.88408126
  when "001011000100"=> s <="111100010100"; -- Argumento 708 Funcion 0.88479710
  when "001011000101"=> s <="111100010101"; -- Argumento 709 Funcion 0.88551086
  when "001011000110"=> s <="111100010110"; -- Argumento 710 Funcion 0.88622253
  when "001011000111"=> s <="111100011000"; -- Argumento 711 Funcion 0.88693212
  when "001011001000"=> s <="111100011001"; -- Argumento 712 Funcion 0.88763962
  when "001011001001"=> s <="111100011011"; -- Argumento 713 Funcion 0.88834503
  when "001011001010"=> s <="111100011100"; -- Argumento 714 Funcion 0.88904836
  when "001011001011"=> s <="111100011110"; -- Argumento 715 Funcion 0.88974959
  when "001011001100"=> s <="111100011111"; -- Argumento 716 Funcion 0.89044872
  when "001011001101"=> s <="111100100001"; -- Argumento 717 Funcion 0.89114576
  when "001011001110"=> s <="111100100010"; -- Argumento 718 Funcion 0.89184071
  when "001011001111"=> s <="111100100011"; -- Argumento 719 Funcion 0.89253356
  when "001011010000"=> s <="111100100101"; -- Argumento 720 Funcion 0.89322430
  when "001011010001"=> s <="111100100110"; -- Argumento 721 Funcion 0.89391295
  when "001011010010"=> s <="111100101000"; -- Argumento 722 Funcion 0.89459949
  when "001011010011"=> s <="111100101001"; -- Argumento 723 Funcion 0.89528392
  when "001011010100"=> s <="111100101010"; -- Argumento 724 Funcion 0.89596625
  when "001011010101"=> s <="111100101100"; -- Argumento 725 Funcion 0.89664647
  when "001011010110"=> s <="111100101101"; -- Argumento 726 Funcion 0.89732458
  when "001011010111"=> s <="111100101111"; -- Argumento 727 Funcion 0.89800058
  when "001011011000"=> s <="111100110000"; -- Argumento 728 Funcion 0.89867447
  when "001011011001"=> s <="111100110001"; -- Argumento 729 Funcion 0.89934624
  when "001011011010"=> s <="111100110011"; -- Argumento 730 Funcion 0.90001589
  when "001011011011"=> s <="111100110100"; -- Argumento 731 Funcion 0.90068343
  when "001011011100"=> s <="111100110101"; -- Argumento 732 Funcion 0.90134885
  when "001011011101"=> s <="111100110111"; -- Argumento 733 Funcion 0.90201214
  when "001011011110"=> s <="111100111000"; -- Argumento 734 Funcion 0.90267332
  when "001011011111"=> s <="111100111010"; -- Argumento 735 Funcion 0.90333237
  when "001011100000"=> s <="111100111011"; -- Argumento 736 Funcion 0.90398929
  when "001011100001"=> s <="111100111100"; -- Argumento 737 Funcion 0.90464409
  when "001011100010"=> s <="111100111110"; -- Argumento 738 Funcion 0.90529676
  when "001011100011"=> s <="111100111111"; -- Argumento 739 Funcion 0.90594730
  when "001011100100"=> s <="111101000000"; -- Argumento 740 Funcion 0.90659570
  when "001011100101"=> s <="111101000010"; -- Argumento 741 Funcion 0.90724198
  when "001011100110"=> s <="111101000011"; -- Argumento 742 Funcion 0.90788612
  when "001011100111"=> s <="111101000100"; -- Argumento 743 Funcion 0.90852812
  when "001011101000"=> s <="111101000101"; -- Argumento 744 Funcion 0.90916798
  when "001011101001"=> s <="111101000111"; -- Argumento 745 Funcion 0.90980571
  when "001011101010"=> s <="111101001000"; -- Argumento 746 Funcion 0.91044129
  when "001011101011"=> s <="111101001001"; -- Argumento 747 Funcion 0.91107473
  when "001011101100"=> s <="111101001011"; -- Argumento 748 Funcion 0.91170603
  when "001011101101"=> s <="111101001100"; -- Argumento 749 Funcion 0.91233518
  when "001011101110"=> s <="111101001101"; -- Argumento 750 Funcion 0.91296219
  when "001011101111"=> s <="111101001111"; -- Argumento 751 Funcion 0.91358705
  when "001011110000"=> s <="111101010000"; -- Argumento 752 Funcion 0.91420976
  when "001011110001"=> s <="111101010001"; -- Argumento 753 Funcion 0.91483031
  when "001011110010"=> s <="111101010010"; -- Argumento 754 Funcion 0.91544872
  when "001011110011"=> s <="111101010100"; -- Argumento 755 Funcion 0.91606497
  when "001011110100"=> s <="111101010101"; -- Argumento 756 Funcion 0.91667906
  when "001011110101"=> s <="111101010110"; -- Argumento 757 Funcion 0.91729100
  when "001011110110"=> s <="111101010111"; -- Argumento 758 Funcion 0.91790078
  when "001011110111"=> s <="111101011001"; -- Argumento 759 Funcion 0.91850839
  when "001011111000"=> s <="111101011010"; -- Argumento 760 Funcion 0.91911385
  when "001011111001"=> s <="111101011011"; -- Argumento 761 Funcion 0.91971715
  when "001011111010"=> s <="111101011100"; -- Argumento 762 Funcion 0.92031828
  when "001011111011"=> s <="111101011110"; -- Argumento 763 Funcion 0.92091724
  when "001011111100"=> s <="111101011111"; -- Argumento 764 Funcion 0.92151404
  when "001011111101"=> s <="111101100000"; -- Argumento 765 Funcion 0.92210867
  when "001011111110"=> s <="111101100001"; -- Argumento 766 Funcion 0.92270113
  when "001011111111"=> s <="111101100010"; -- Argumento 767 Funcion 0.92329142
  when "001100000000"=> s <="111101100100"; -- Argumento 768 Funcion 0.92387953
  when "001100000001"=> s <="111101100101"; -- Argumento 769 Funcion 0.92446547
  when "001100000010"=> s <="111101100110"; -- Argumento 770 Funcion 0.92504924
  when "001100000011"=> s <="111101100111"; -- Argumento 771 Funcion 0.92563083
  when "001100000100"=> s <="111101101000"; -- Argumento 772 Funcion 0.92621024
  when "001100000101"=> s <="111101101010"; -- Argumento 773 Funcion 0.92678747
  when "001100000110"=> s <="111101101011"; -- Argumento 774 Funcion 0.92736253
  when "001100000111"=> s <="111101101100"; -- Argumento 775 Funcion 0.92793539
  when "001100001000"=> s <="111101101101"; -- Argumento 776 Funcion 0.92850608
  when "001100001001"=> s <="111101101110"; -- Argumento 777 Funcion 0.92907458
  when "001100001010"=> s <="111101101111"; -- Argumento 778 Funcion 0.92964090
  when "001100001011"=> s <="111101110001"; -- Argumento 779 Funcion 0.93020502
  when "001100001100"=> s <="111101110010"; -- Argumento 780 Funcion 0.93076696
  when "001100001101"=> s <="111101110011"; -- Argumento 781 Funcion 0.93132671
  when "001100001110"=> s <="111101110100"; -- Argumento 782 Funcion 0.93188427
  when "001100001111"=> s <="111101110101"; -- Argumento 783 Funcion 0.93243963
  when "001100010000"=> s <="111101110110"; -- Argumento 784 Funcion 0.93299280
  when "001100010001"=> s <="111101110111"; -- Argumento 785 Funcion 0.93354377
  when "001100010010"=> s <="111101111001"; -- Argumento 786 Funcion 0.93409255
  when "001100010011"=> s <="111101111010"; -- Argumento 787 Funcion 0.93463913
  when "001100010100"=> s <="111101111011"; -- Argumento 788 Funcion 0.93518351
  when "001100010101"=> s <="111101111100"; -- Argumento 789 Funcion 0.93572569
  when "001100010110"=> s <="111101111101"; -- Argumento 790 Funcion 0.93626567
  when "001100010111"=> s <="111101111110"; -- Argumento 791 Funcion 0.93680344
  when "001100011000"=> s <="111101111111"; -- Argumento 792 Funcion 0.93733901
  when "001100011001"=> s <="111110000000"; -- Argumento 793 Funcion 0.93787238
  when "001100011010"=> s <="111110000001"; -- Argumento 794 Funcion 0.93840353
  when "001100011011"=> s <="111110000010"; -- Argumento 795 Funcion 0.93893248
  when "001100011100"=> s <="111110000100"; -- Argumento 796 Funcion 0.93945922
  when "001100011101"=> s <="111110000101"; -- Argumento 797 Funcion 0.93998375
  when "001100011110"=> s <="111110000110"; -- Argumento 798 Funcion 0.94050607
  when "001100011111"=> s <="111110000111"; -- Argumento 799 Funcion 0.94102618
  when "001100100000"=> s <="111110001000"; -- Argumento 800 Funcion 0.94154407
  when "001100100001"=> s <="111110001001"; -- Argumento 801 Funcion 0.94205974
  when "001100100010"=> s <="111110001010"; -- Argumento 802 Funcion 0.94257320
  when "001100100011"=> s <="111110001011"; -- Argumento 803 Funcion 0.94308444
  when "001100100100"=> s <="111110001100"; -- Argumento 804 Funcion 0.94359346
  when "001100100101"=> s <="111110001101"; -- Argumento 805 Funcion 0.94410026
  when "001100100110"=> s <="111110001110"; -- Argumento 806 Funcion 0.94460484
  when "001100100111"=> s <="111110001111"; -- Argumento 807 Funcion 0.94510719
  when "001100101000"=> s <="111110010000"; -- Argumento 808 Funcion 0.94560733
  when "001100101001"=> s <="111110010001"; -- Argumento 809 Funcion 0.94610523
  when "001100101010"=> s <="111110010010"; -- Argumento 810 Funcion 0.94660091
  when "001100101011"=> s <="111110010011"; -- Argumento 811 Funcion 0.94709437
  when "001100101100"=> s <="111110010100"; -- Argumento 812 Funcion 0.94758559
  when "001100101101"=> s <="111110010101"; -- Argumento 813 Funcion 0.94807459
  when "001100101110"=> s <="111110010110"; -- Argumento 814 Funcion 0.94856135
  when "001100101111"=> s <="111110010111"; -- Argumento 815 Funcion 0.94904588
  when "001100110000"=> s <="111110011000"; -- Argumento 816 Funcion 0.94952818
  when "001100110001"=> s <="111110011001"; -- Argumento 817 Funcion 0.95000825
  when "001100110010"=> s <="111110011010"; -- Argumento 818 Funcion 0.95048607
  when "001100110011"=> s <="111110011011"; -- Argumento 819 Funcion 0.95096167
  when "001100110100"=> s <="111110011100"; -- Argumento 820 Funcion 0.95143502
  when "001100110101"=> s <="111110011101"; -- Argumento 821 Funcion 0.95190614
  when "001100110110"=> s <="111110011110"; -- Argumento 822 Funcion 0.95237501
  when "001100110111"=> s <="111110011111"; -- Argumento 823 Funcion 0.95284165
  when "001100111000"=> s <="111110100000"; -- Argumento 824 Funcion 0.95330604
  when "001100111001"=> s <="111110100001"; -- Argumento 825 Funcion 0.95376819
  when "001100111010"=> s <="111110100010"; -- Argumento 826 Funcion 0.95422810
  when "001100111011"=> s <="111110100011"; -- Argumento 827 Funcion 0.95468575
  when "001100111100"=> s <="111110100100"; -- Argumento 828 Funcion 0.95514117
  when "001100111101"=> s <="111110100101"; -- Argumento 829 Funcion 0.95559433
  when "001100111110"=> s <="111110100101"; -- Argumento 830 Funcion 0.95604525
  when "001100111111"=> s <="111110100110"; -- Argumento 831 Funcion 0.95649392
  when "001101000000"=> s <="111110100111"; -- Argumento 832 Funcion 0.95694034
  when "001101000001"=> s <="111110101000"; -- Argumento 833 Funcion 0.95738450
  when "001101000010"=> s <="111110101001"; -- Argumento 834 Funcion 0.95782641
  when "001101000011"=> s <="111110101010"; -- Argumento 835 Funcion 0.95826607
  when "001101000100"=> s <="111110101011"; -- Argumento 836 Funcion 0.95870347
  when "001101000101"=> s <="111110101100"; -- Argumento 837 Funcion 0.95913862
  when "001101000110"=> s <="111110101101"; -- Argumento 838 Funcion 0.95957151
  when "001101000111"=> s <="111110101110"; -- Argumento 839 Funcion 0.96000215
  when "001101001000"=> s <="111110101110"; -- Argumento 840 Funcion 0.96043052
  when "001101001001"=> s <="111110101111"; -- Argumento 841 Funcion 0.96085663
  when "001101001010"=> s <="111110110000"; -- Argumento 842 Funcion 0.96128049
  when "001101001011"=> s <="111110110001"; -- Argumento 843 Funcion 0.96170208
  when "001101001100"=> s <="111110110010"; -- Argumento 844 Funcion 0.96212140
  when "001101001101"=> s <="111110110011"; -- Argumento 845 Funcion 0.96253847
  when "001101001110"=> s <="111110110100"; -- Argumento 846 Funcion 0.96295327
  when "001101001111"=> s <="111110110100"; -- Argumento 847 Funcion 0.96336580
  when "001101010000"=> s <="111110110101"; -- Argumento 848 Funcion 0.96377607
  when "001101010001"=> s <="111110110110"; -- Argumento 849 Funcion 0.96418406
  when "001101010010"=> s <="111110110111"; -- Argumento 850 Funcion 0.96458979
  when "001101010011"=> s <="111110111000"; -- Argumento 851 Funcion 0.96499325
  when "001101010100"=> s <="111110111001"; -- Argumento 852 Funcion 0.96539444
  when "001101010101"=> s <="111110111001"; -- Argumento 853 Funcion 0.96579336
  when "001101010110"=> s <="111110111010"; -- Argumento 854 Funcion 0.96619000
  when "001101010111"=> s <="111110111011"; -- Argumento 855 Funcion 0.96658437
  when "001101011000"=> s <="111110111100"; -- Argumento 856 Funcion 0.96697647
  when "001101011001"=> s <="111110111101"; -- Argumento 857 Funcion 0.96736629
  when "001101011010"=> s <="111110111101"; -- Argumento 858 Funcion 0.96775384
  when "001101011011"=> s <="111110111110"; -- Argumento 859 Funcion 0.96813910
  when "001101011100"=> s <="111110111111"; -- Argumento 860 Funcion 0.96852209
  when "001101011101"=> s <="111111000000"; -- Argumento 861 Funcion 0.96890280
  when "001101011110"=> s <="111111000001"; -- Argumento 862 Funcion 0.96928124
  when "001101011111"=> s <="111111000001"; -- Argumento 863 Funcion 0.96965739
  when "001101100000"=> s <="111111000010"; -- Argumento 864 Funcion 0.97003125
  when "001101100001"=> s <="111111000011"; -- Argumento 865 Funcion 0.97040284
  when "001101100010"=> s <="111111000100"; -- Argumento 866 Funcion 0.97077214
  when "001101100011"=> s <="111111000100"; -- Argumento 867 Funcion 0.97113916
  when "001101100100"=> s <="111111000101"; -- Argumento 868 Funcion 0.97150389
  when "001101100101"=> s <="111111000110"; -- Argumento 869 Funcion 0.97186634
  when "001101100110"=> s <="111111000111"; -- Argumento 870 Funcion 0.97222650
  when "001101100111"=> s <="111111000111"; -- Argumento 871 Funcion 0.97258437
  when "001101101000"=> s <="111111001000"; -- Argumento 872 Funcion 0.97293995
  when "001101101001"=> s <="111111001001"; -- Argumento 873 Funcion 0.97329325
  when "001101101010"=> s <="111111001010"; -- Argumento 874 Funcion 0.97364425
  when "001101101011"=> s <="111111001010"; -- Argumento 875 Funcion 0.97399296
  when "001101101100"=> s <="111111001011"; -- Argumento 876 Funcion 0.97433938
  when "001101101101"=> s <="111111001100"; -- Argumento 877 Funcion 0.97468351
  when "001101101110"=> s <="111111001100"; -- Argumento 878 Funcion 0.97502535
  when "001101101111"=> s <="111111001101"; -- Argumento 879 Funcion 0.97536489
  when "001101110000"=> s <="111111001110"; -- Argumento 880 Funcion 0.97570213
  when "001101110001"=> s <="111111001110"; -- Argumento 881 Funcion 0.97603708
  when "001101110010"=> s <="111111001111"; -- Argumento 882 Funcion 0.97636973
  when "001101110011"=> s <="111111010000"; -- Argumento 883 Funcion 0.97670009
  when "001101110100"=> s <="111111010000"; -- Argumento 884 Funcion 0.97702814
  when "001101110101"=> s <="111111010001"; -- Argumento 885 Funcion 0.97735390
  when "001101110110"=> s <="111111010010"; -- Argumento 886 Funcion 0.97767736
  when "001101110111"=> s <="111111010010"; -- Argumento 887 Funcion 0.97799851
  when "001101111000"=> s <="111111010011"; -- Argumento 888 Funcion 0.97831737
  when "001101111001"=> s <="111111010100"; -- Argumento 889 Funcion 0.97863392
  when "001101111010"=> s <="111111010100"; -- Argumento 890 Funcion 0.97894818
  when "001101111011"=> s <="111111010101"; -- Argumento 891 Funcion 0.97926012
  when "001101111100"=> s <="111111010110"; -- Argumento 892 Funcion 0.97956977
  when "001101111101"=> s <="111111010110"; -- Argumento 893 Funcion 0.97987710
  when "001101111110"=> s <="111111010111"; -- Argumento 894 Funcion 0.98018214
  when "001101111111"=> s <="111111011000"; -- Argumento 895 Funcion 0.98048486
  when "001110000000"=> s <="111111011000"; -- Argumento 896 Funcion 0.98078528
  when "001110000001"=> s <="111111011001"; -- Argumento 897 Funcion 0.98108339
  when "001110000010"=> s <="111111011001"; -- Argumento 898 Funcion 0.98137919
  when "001110000011"=> s <="111111011010"; -- Argumento 899 Funcion 0.98167269
  when "001110000100"=> s <="111111011011"; -- Argumento 900 Funcion 0.98196387
  when "001110000101"=> s <="111111011011"; -- Argumento 901 Funcion 0.98225274
  when "001110000110"=> s <="111111011100"; -- Argumento 902 Funcion 0.98253930
  when "001110000111"=> s <="111111011100"; -- Argumento 903 Funcion 0.98282355
  when "001110001000"=> s <="111111011101"; -- Argumento 904 Funcion 0.98310549
  when "001110001001"=> s <="111111011101"; -- Argumento 905 Funcion 0.98338511
  when "001110001010"=> s <="111111011110"; -- Argumento 906 Funcion 0.98366242
  when "001110001011"=> s <="111111011111"; -- Argumento 907 Funcion 0.98393741
  when "001110001100"=> s <="111111011111"; -- Argumento 908 Funcion 0.98421009
  when "001110001101"=> s <="111111100000"; -- Argumento 909 Funcion 0.98448046
  when "001110001110"=> s <="111111100000"; -- Argumento 910 Funcion 0.98474850
  when "001110001111"=> s <="111111100001"; -- Argumento 911 Funcion 0.98501423
  when "001110010000"=> s <="111111100001"; -- Argumento 912 Funcion 0.98527764
  when "001110010001"=> s <="111111100010"; -- Argumento 913 Funcion 0.98553874
  when "001110010010"=> s <="111111100010"; -- Argumento 914 Funcion 0.98579751
  when "001110010011"=> s <="111111100011"; -- Argumento 915 Funcion 0.98605396
  when "001110010100"=> s <="111111100011"; -- Argumento 916 Funcion 0.98630810
  when "001110010101"=> s <="111111100100"; -- Argumento 917 Funcion 0.98655991
  when "001110010110"=> s <="111111100100"; -- Argumento 918 Funcion 0.98680940
  when "001110010111"=> s <="111111100101"; -- Argumento 919 Funcion 0.98705657
  when "001110011000"=> s <="111111100101"; -- Argumento 920 Funcion 0.98730142
  when "001110011001"=> s <="111111100110"; -- Argumento 921 Funcion 0.98754394
  when "001110011010"=> s <="111111100110"; -- Argumento 922 Funcion 0.98778414
  when "001110011011"=> s <="111111100111"; -- Argumento 923 Funcion 0.98802202
  when "001110011100"=> s <="111111100111"; -- Argumento 924 Funcion 0.98825757
  when "001110011101"=> s <="111111101000"; -- Argumento 925 Funcion 0.98849079
  when "001110011110"=> s <="111111101000"; -- Argumento 926 Funcion 0.98872169
  when "001110011111"=> s <="111111101001"; -- Argumento 927 Funcion 0.98895026
  when "001110100000"=> s <="111111101001"; -- Argumento 928 Funcion 0.98917651
  when "001110100001"=> s <="111111101010"; -- Argumento 929 Funcion 0.98940043
  when "001110100010"=> s <="111111101010"; -- Argumento 930 Funcion 0.98962202
  when "001110100011"=> s <="111111101011"; -- Argumento 931 Funcion 0.98984128
  when "001110100100"=> s <="111111101011"; -- Argumento 932 Funcion 0.99005821
  when "001110100101"=> s <="111111101100"; -- Argumento 933 Funcion 0.99027281
  when "001110100110"=> s <="111111101100"; -- Argumento 934 Funcion 0.99048508
  when "001110100111"=> s <="111111101100"; -- Argumento 935 Funcion 0.99069503
  when "001110101000"=> s <="111111101101"; -- Argumento 936 Funcion 0.99090264
  when "001110101001"=> s <="111111101101"; -- Argumento 937 Funcion 0.99110791
  when "001110101010"=> s <="111111101110"; -- Argumento 938 Funcion 0.99131086
  when "001110101011"=> s <="111111101110"; -- Argumento 939 Funcion 0.99151147
  when "001110101100"=> s <="111111101111"; -- Argumento 940 Funcion 0.99170975
  when "001110101101"=> s <="111111101111"; -- Argumento 941 Funcion 0.99190570
  when "001110101110"=> s <="111111101111"; -- Argumento 942 Funcion 0.99209931
  when "001110101111"=> s <="111111110000"; -- Argumento 943 Funcion 0.99229059
  when "001110110000"=> s <="111111110000"; -- Argumento 944 Funcion 0.99247953
  when "001110110001"=> s <="111111110000"; -- Argumento 945 Funcion 0.99266614
  when "001110110010"=> s <="111111110001"; -- Argumento 946 Funcion 0.99285041
  when "001110110011"=> s <="111111110001"; -- Argumento 947 Funcion 0.99303235
  when "001110110100"=> s <="111111110010"; -- Argumento 948 Funcion 0.99321195
  when "001110110101"=> s <="111111110010"; -- Argumento 949 Funcion 0.99338921
  when "001110110110"=> s <="111111110010"; -- Argumento 950 Funcion 0.99356414
  when "001110110111"=> s <="111111110011"; -- Argumento 951 Funcion 0.99373672
  when "001110111000"=> s <="111111110011"; -- Argumento 952 Funcion 0.99390697
  when "001110111001"=> s <="111111110011"; -- Argumento 953 Funcion 0.99407488
  when "001110111010"=> s <="111111110100"; -- Argumento 954 Funcion 0.99424045
  when "001110111011"=> s <="111111110100"; -- Argumento 955 Funcion 0.99440368
  when "001110111100"=> s <="111111110100"; -- Argumento 956 Funcion 0.99456457
  when "001110111101"=> s <="111111110101"; -- Argumento 957 Funcion 0.99472312
  when "001110111110"=> s <="111111110101"; -- Argumento 958 Funcion 0.99487933
  when "001110111111"=> s <="111111110101"; -- Argumento 959 Funcion 0.99503320
  when "001111000000"=> s <="111111110110"; -- Argumento 960 Funcion 0.99518473
  when "001111000001"=> s <="111111110110"; -- Argumento 961 Funcion 0.99533391
  when "001111000010"=> s <="111111110110"; -- Argumento 962 Funcion 0.99548076
  when "001111000011"=> s <="111111110111"; -- Argumento 963 Funcion 0.99562526
  when "001111000100"=> s <="111111110111"; -- Argumento 964 Funcion 0.99576741
  when "001111000101"=> s <="111111110111"; -- Argumento 965 Funcion 0.99590723
  when "001111000110"=> s <="111111110111"; -- Argumento 966 Funcion 0.99604470
  when "001111000111"=> s <="111111111000"; -- Argumento 967 Funcion 0.99617983
  when "001111001000"=> s <="111111111000"; -- Argumento 968 Funcion 0.99631261
  when "001111001001"=> s <="111111111000"; -- Argumento 969 Funcion 0.99644305
  when "001111001010"=> s <="111111111000"; -- Argumento 970 Funcion 0.99657115
  when "001111001011"=> s <="111111111001"; -- Argumento 971 Funcion 0.99669690
  when "001111001100"=> s <="111111111001"; -- Argumento 972 Funcion 0.99682030
  when "001111001101"=> s <="111111111001"; -- Argumento 973 Funcion 0.99694136
  when "001111001110"=> s <="111111111001"; -- Argumento 974 Funcion 0.99706007
  when "001111001111"=> s <="111111111010"; -- Argumento 975 Funcion 0.99717644
  when "001111010000"=> s <="111111111010"; -- Argumento 976 Funcion 0.99729046
  when "001111010001"=> s <="111111111010"; -- Argumento 977 Funcion 0.99740213
  when "001111010010"=> s <="111111111010"; -- Argumento 978 Funcion 0.99751146
  when "001111010011"=> s <="111111111011"; -- Argumento 979 Funcion 0.99761844
  when "001111010100"=> s <="111111111011"; -- Argumento 980 Funcion 0.99772307
  when "001111010101"=> s <="111111111011"; -- Argumento 981 Funcion 0.99782535
  when "001111010110"=> s <="111111111011"; -- Argumento 982 Funcion 0.99792529
  when "001111010111"=> s <="111111111011"; -- Argumento 983 Funcion 0.99802287
  when "001111011000"=> s <="111111111100"; -- Argumento 984 Funcion 0.99811811
  when "001111011001"=> s <="111111111100"; -- Argumento 985 Funcion 0.99821100
  when "001111011010"=> s <="111111111100"; -- Argumento 986 Funcion 0.99830154
  when "001111011011"=> s <="111111111100"; -- Argumento 987 Funcion 0.99838974
  when "001111011100"=> s <="111111111100"; -- Argumento 988 Funcion 0.99847558
  when "001111011101"=> s <="111111111101"; -- Argumento 989 Funcion 0.99855907
  when "001111011110"=> s <="111111111101"; -- Argumento 990 Funcion 0.99864022
  when "001111011111"=> s <="111111111101"; -- Argumento 991 Funcion 0.99871901
  when "001111100000"=> s <="111111111101"; -- Argumento 992 Funcion 0.99879546
  when "001111100001"=> s <="111111111101"; -- Argumento 993 Funcion 0.99886955
  when "001111100010"=> s <="111111111101"; -- Argumento 994 Funcion 0.99894129
  when "001111100011"=> s <="111111111101"; -- Argumento 995 Funcion 0.99901069
  when "001111100100"=> s <="111111111110"; -- Argumento 996 Funcion 0.99907773
  when "001111100101"=> s <="111111111110"; -- Argumento 997 Funcion 0.99914242
  when "001111100110"=> s <="111111111110"; -- Argumento 998 Funcion 0.99920476
  when "001111100111"=> s <="111111111110"; -- Argumento 999 Funcion 0.99926475
  when "001111101000"=> s <="111111111110"; -- Argumento 1000 Funcion 0.99932238
  when "001111101001"=> s <="111111111110"; -- Argumento 1001 Funcion 0.99937767
  when "001111101010"=> s <="111111111110"; -- Argumento 1002 Funcion 0.99943060
  when "001111101011"=> s <="111111111110"; -- Argumento 1003 Funcion 0.99948119
  when "001111101100"=> s <="111111111111"; -- Argumento 1004 Funcion 0.99952942
  when "001111101101"=> s <="111111111111"; -- Argumento 1005 Funcion 0.99957530
  when "001111101110"=> s <="111111111111"; -- Argumento 1006 Funcion 0.99961882
  when "001111101111"=> s <="111111111111"; -- Argumento 1007 Funcion 0.99966000
  when "001111110000"=> s <="111111111111"; -- Argumento 1008 Funcion 0.99969882
  when "001111110001"=> s <="111111111111"; -- Argumento 1009 Funcion 0.99973529
  when "001111110010"=> s <="111111111111"; -- Argumento 1010 Funcion 0.99976941
  when "001111110011"=> s <="111111111111"; -- Argumento 1011 Funcion 0.99980117
  when "001111110100"=> s <="111111111111"; -- Argumento 1012 Funcion 0.99983058
  when "001111110101"=> s <="111111111111"; -- Argumento 1013 Funcion 0.99985764
  when "001111110110"=> s <="111111111111"; -- Argumento 1014 Funcion 0.99988235
  when "001111110111"=> s <="111111111111"; -- Argumento 1015 Funcion 0.99990470
  when "001111111000"=> s <="111111111111"; -- Argumento 1016 Funcion 0.99992470
  when "001111111001"=> s <="111111111111"; -- Argumento 1017 Funcion 0.99994235
  when "001111111010"=> s <="111111111111"; -- Argumento 1018 Funcion 0.99995764
  when "001111111011"=> s <="111111111111"; -- Argumento 1019 Funcion 0.99997059
  when "001111111100"=> s <="111111111111"; -- Argumento 1020 Funcion 0.99998118
  when "001111111101"=> s <="111111111111"; -- Argumento 1021 Funcion 0.99998941
  when "001111111110"=> s <="111111111111"; -- Argumento 1022 Funcion 0.99999529
  when "001111111111"=> s <="111111111111"; -- Argumento 1023 Funcion 0.99999882
  when "010000000000"=> s <="111111111111"; -- Argumento 1024 Funcion 1.00000000
  when "010000000001"=> s <="111111111111"; -- Argumento 1025 Funcion 0.99999882
  when "010000000010"=> s <="111111111111"; -- Argumento 1026 Funcion 0.99999529
  when "010000000011"=> s <="111111111111"; -- Argumento 1027 Funcion 0.99998941
  when "010000000100"=> s <="111111111111"; -- Argumento 1028 Funcion 0.99998118
  when "010000000101"=> s <="111111111111"; -- Argumento 1029 Funcion 0.99997059
  when "010000000110"=> s <="111111111111"; -- Argumento 1030 Funcion 0.99995764
  when "010000000111"=> s <="111111111111"; -- Argumento 1031 Funcion 0.99994235
  when "010000001000"=> s <="111111111111"; -- Argumento 1032 Funcion 0.99992470
  when "010000001001"=> s <="111111111111"; -- Argumento 1033 Funcion 0.99990470
  when "010000001010"=> s <="111111111111"; -- Argumento 1034 Funcion 0.99988235
  when "010000001011"=> s <="111111111111"; -- Argumento 1035 Funcion 0.99985764
  when "010000001100"=> s <="111111111111"; -- Argumento 1036 Funcion 0.99983058
  when "010000001101"=> s <="111111111111"; -- Argumento 1037 Funcion 0.99980117
  when "010000001110"=> s <="111111111111"; -- Argumento 1038 Funcion 0.99976941
  when "010000001111"=> s <="111111111111"; -- Argumento 1039 Funcion 0.99973529
  when "010000010000"=> s <="111111111111"; -- Argumento 1040 Funcion 0.99969882
  when "010000010001"=> s <="111111111111"; -- Argumento 1041 Funcion 0.99966000
  when "010000010010"=> s <="111111111111"; -- Argumento 1042 Funcion 0.99961882
  when "010000010011"=> s <="111111111111"; -- Argumento 1043 Funcion 0.99957530
  when "010000010100"=> s <="111111111111"; -- Argumento 1044 Funcion 0.99952942
  when "010000010101"=> s <="111111111110"; -- Argumento 1045 Funcion 0.99948119
  when "010000010110"=> s <="111111111110"; -- Argumento 1046 Funcion 0.99943060
  when "010000010111"=> s <="111111111110"; -- Argumento 1047 Funcion 0.99937767
  when "010000011000"=> s <="111111111110"; -- Argumento 1048 Funcion 0.99932238
  when "010000011001"=> s <="111111111110"; -- Argumento 1049 Funcion 0.99926475
  when "010000011010"=> s <="111111111110"; -- Argumento 1050 Funcion 0.99920476
  when "010000011011"=> s <="111111111110"; -- Argumento 1051 Funcion 0.99914242
  when "010000011100"=> s <="111111111110"; -- Argumento 1052 Funcion 0.99907773
  when "010000011101"=> s <="111111111101"; -- Argumento 1053 Funcion 0.99901069
  when "010000011110"=> s <="111111111101"; -- Argumento 1054 Funcion 0.99894129
  when "010000011111"=> s <="111111111101"; -- Argumento 1055 Funcion 0.99886955
  when "010000100000"=> s <="111111111101"; -- Argumento 1056 Funcion 0.99879546
  when "010000100001"=> s <="111111111101"; -- Argumento 1057 Funcion 0.99871901
  when "010000100010"=> s <="111111111101"; -- Argumento 1058 Funcion 0.99864022
  when "010000100011"=> s <="111111111101"; -- Argumento 1059 Funcion 0.99855907
  when "010000100100"=> s <="111111111100"; -- Argumento 1060 Funcion 0.99847558
  when "010000100101"=> s <="111111111100"; -- Argumento 1061 Funcion 0.99838974
  when "010000100110"=> s <="111111111100"; -- Argumento 1062 Funcion 0.99830154
  when "010000100111"=> s <="111111111100"; -- Argumento 1063 Funcion 0.99821100
  when "010000101000"=> s <="111111111100"; -- Argumento 1064 Funcion 0.99811811
  when "010000101001"=> s <="111111111011"; -- Argumento 1065 Funcion 0.99802287
  when "010000101010"=> s <="111111111011"; -- Argumento 1066 Funcion 0.99792529
  when "010000101011"=> s <="111111111011"; -- Argumento 1067 Funcion 0.99782535
  when "010000101100"=> s <="111111111011"; -- Argumento 1068 Funcion 0.99772307
  when "010000101101"=> s <="111111111011"; -- Argumento 1069 Funcion 0.99761844
  when "010000101110"=> s <="111111111010"; -- Argumento 1070 Funcion 0.99751146
  when "010000101111"=> s <="111111111010"; -- Argumento 1071 Funcion 0.99740213
  when "010000110000"=> s <="111111111010"; -- Argumento 1072 Funcion 0.99729046
  when "010000110001"=> s <="111111111010"; -- Argumento 1073 Funcion 0.99717644
  when "010000110010"=> s <="111111111001"; -- Argumento 1074 Funcion 0.99706007
  when "010000110011"=> s <="111111111001"; -- Argumento 1075 Funcion 0.99694136
  when "010000110100"=> s <="111111111001"; -- Argumento 1076 Funcion 0.99682030
  when "010000110101"=> s <="111111111001"; -- Argumento 1077 Funcion 0.99669690
  when "010000110110"=> s <="111111111000"; -- Argumento 1078 Funcion 0.99657115
  when "010000110111"=> s <="111111111000"; -- Argumento 1079 Funcion 0.99644305
  when "010000111000"=> s <="111111111000"; -- Argumento 1080 Funcion 0.99631261
  when "010000111001"=> s <="111111111000"; -- Argumento 1081 Funcion 0.99617983
  when "010000111010"=> s <="111111110111"; -- Argumento 1082 Funcion 0.99604470
  when "010000111011"=> s <="111111110111"; -- Argumento 1083 Funcion 0.99590723
  when "010000111100"=> s <="111111110111"; -- Argumento 1084 Funcion 0.99576741
  when "010000111101"=> s <="111111110111"; -- Argumento 1085 Funcion 0.99562526
  when "010000111110"=> s <="111111110110"; -- Argumento 1086 Funcion 0.99548076
  when "010000111111"=> s <="111111110110"; -- Argumento 1087 Funcion 0.99533391
  when "010001000000"=> s <="111111110110"; -- Argumento 1088 Funcion 0.99518473
  when "010001000001"=> s <="111111110101"; -- Argumento 1089 Funcion 0.99503320
  when "010001000010"=> s <="111111110101"; -- Argumento 1090 Funcion 0.99487933
  when "010001000011"=> s <="111111110101"; -- Argumento 1091 Funcion 0.99472312
  when "010001000100"=> s <="111111110100"; -- Argumento 1092 Funcion 0.99456457
  when "010001000101"=> s <="111111110100"; -- Argumento 1093 Funcion 0.99440368
  when "010001000110"=> s <="111111110100"; -- Argumento 1094 Funcion 0.99424045
  when "010001000111"=> s <="111111110011"; -- Argumento 1095 Funcion 0.99407488
  when "010001001000"=> s <="111111110011"; -- Argumento 1096 Funcion 0.99390697
  when "010001001001"=> s <="111111110011"; -- Argumento 1097 Funcion 0.99373672
  when "010001001010"=> s <="111111110010"; -- Argumento 1098 Funcion 0.99356414
  when "010001001011"=> s <="111111110010"; -- Argumento 1099 Funcion 0.99338921
  when "010001001100"=> s <="111111110010"; -- Argumento 1100 Funcion 0.99321195
  when "010001001101"=> s <="111111110001"; -- Argumento 1101 Funcion 0.99303235
  when "010001001110"=> s <="111111110001"; -- Argumento 1102 Funcion 0.99285041
  when "010001001111"=> s <="111111110000"; -- Argumento 1103 Funcion 0.99266614
  when "010001010000"=> s <="111111110000"; -- Argumento 1104 Funcion 0.99247953
  when "010001010001"=> s <="111111110000"; -- Argumento 1105 Funcion 0.99229059
  when "010001010010"=> s <="111111101111"; -- Argumento 1106 Funcion 0.99209931
  when "010001010011"=> s <="111111101111"; -- Argumento 1107 Funcion 0.99190570
  when "010001010100"=> s <="111111101111"; -- Argumento 1108 Funcion 0.99170975
  when "010001010101"=> s <="111111101110"; -- Argumento 1109 Funcion 0.99151147
  when "010001010110"=> s <="111111101110"; -- Argumento 1110 Funcion 0.99131086
  when "010001010111"=> s <="111111101101"; -- Argumento 1111 Funcion 0.99110791
  when "010001011000"=> s <="111111101101"; -- Argumento 1112 Funcion 0.99090264
  when "010001011001"=> s <="111111101100"; -- Argumento 1113 Funcion 0.99069503
  when "010001011010"=> s <="111111101100"; -- Argumento 1114 Funcion 0.99048508
  when "010001011011"=> s <="111111101100"; -- Argumento 1115 Funcion 0.99027281
  when "010001011100"=> s <="111111101011"; -- Argumento 1116 Funcion 0.99005821
  when "010001011101"=> s <="111111101011"; -- Argumento 1117 Funcion 0.98984128
  when "010001011110"=> s <="111111101010"; -- Argumento 1118 Funcion 0.98962202
  when "010001011111"=> s <="111111101010"; -- Argumento 1119 Funcion 0.98940043
  when "010001100000"=> s <="111111101001"; -- Argumento 1120 Funcion 0.98917651
  when "010001100001"=> s <="111111101001"; -- Argumento 1121 Funcion 0.98895026
  when "010001100010"=> s <="111111101000"; -- Argumento 1122 Funcion 0.98872169
  when "010001100011"=> s <="111111101000"; -- Argumento 1123 Funcion 0.98849079
  when "010001100100"=> s <="111111100111"; -- Argumento 1124 Funcion 0.98825757
  when "010001100101"=> s <="111111100111"; -- Argumento 1125 Funcion 0.98802202
  when "010001100110"=> s <="111111100110"; -- Argumento 1126 Funcion 0.98778414
  when "010001100111"=> s <="111111100110"; -- Argumento 1127 Funcion 0.98754394
  when "010001101000"=> s <="111111100101"; -- Argumento 1128 Funcion 0.98730142
  when "010001101001"=> s <="111111100101"; -- Argumento 1129 Funcion 0.98705657
  when "010001101010"=> s <="111111100100"; -- Argumento 1130 Funcion 0.98680940
  when "010001101011"=> s <="111111100100"; -- Argumento 1131 Funcion 0.98655991
  when "010001101100"=> s <="111111100011"; -- Argumento 1132 Funcion 0.98630810
  when "010001101101"=> s <="111111100011"; -- Argumento 1133 Funcion 0.98605396
  when "010001101110"=> s <="111111100010"; -- Argumento 1134 Funcion 0.98579751
  when "010001101111"=> s <="111111100010"; -- Argumento 1135 Funcion 0.98553874
  when "010001110000"=> s <="111111100001"; -- Argumento 1136 Funcion 0.98527764
  when "010001110001"=> s <="111111100001"; -- Argumento 1137 Funcion 0.98501423
  when "010001110010"=> s <="111111100000"; -- Argumento 1138 Funcion 0.98474850
  when "010001110011"=> s <="111111100000"; -- Argumento 1139 Funcion 0.98448046
  when "010001110100"=> s <="111111011111"; -- Argumento 1140 Funcion 0.98421009
  when "010001110101"=> s <="111111011111"; -- Argumento 1141 Funcion 0.98393741
  when "010001110110"=> s <="111111011110"; -- Argumento 1142 Funcion 0.98366242
  when "010001110111"=> s <="111111011101"; -- Argumento 1143 Funcion 0.98338511
  when "010001111000"=> s <="111111011101"; -- Argumento 1144 Funcion 0.98310549
  when "010001111001"=> s <="111111011100"; -- Argumento 1145 Funcion 0.98282355
  when "010001111010"=> s <="111111011100"; -- Argumento 1146 Funcion 0.98253930
  when "010001111011"=> s <="111111011011"; -- Argumento 1147 Funcion 0.98225274
  when "010001111100"=> s <="111111011011"; -- Argumento 1148 Funcion 0.98196387
  when "010001111101"=> s <="111111011010"; -- Argumento 1149 Funcion 0.98167269
  when "010001111110"=> s <="111111011001"; -- Argumento 1150 Funcion 0.98137919
  when "010001111111"=> s <="111111011001"; -- Argumento 1151 Funcion 0.98108339
  when "010010000000"=> s <="111111011000"; -- Argumento 1152 Funcion 0.98078528
  when "010010000001"=> s <="111111011000"; -- Argumento 1153 Funcion 0.98048486
  when "010010000010"=> s <="111111010111"; -- Argumento 1154 Funcion 0.98018214
  when "010010000011"=> s <="111111010110"; -- Argumento 1155 Funcion 0.97987710
  when "010010000100"=> s <="111111010110"; -- Argumento 1156 Funcion 0.97956977
  when "010010000101"=> s <="111111010101"; -- Argumento 1157 Funcion 0.97926012
  when "010010000110"=> s <="111111010100"; -- Argumento 1158 Funcion 0.97894818
  when "010010000111"=> s <="111111010100"; -- Argumento 1159 Funcion 0.97863392
  when "010010001000"=> s <="111111010011"; -- Argumento 1160 Funcion 0.97831737
  when "010010001001"=> s <="111111010010"; -- Argumento 1161 Funcion 0.97799851
  when "010010001010"=> s <="111111010010"; -- Argumento 1162 Funcion 0.97767736
  when "010010001011"=> s <="111111010001"; -- Argumento 1163 Funcion 0.97735390
  when "010010001100"=> s <="111111010000"; -- Argumento 1164 Funcion 0.97702814
  when "010010001101"=> s <="111111010000"; -- Argumento 1165 Funcion 0.97670009
  when "010010001110"=> s <="111111001111"; -- Argumento 1166 Funcion 0.97636973
  when "010010001111"=> s <="111111001110"; -- Argumento 1167 Funcion 0.97603708
  when "010010010000"=> s <="111111001110"; -- Argumento 1168 Funcion 0.97570213
  when "010010010001"=> s <="111111001101"; -- Argumento 1169 Funcion 0.97536489
  when "010010010010"=> s <="111111001100"; -- Argumento 1170 Funcion 0.97502535
  when "010010010011"=> s <="111111001100"; -- Argumento 1171 Funcion 0.97468351
  when "010010010100"=> s <="111111001011"; -- Argumento 1172 Funcion 0.97433938
  when "010010010101"=> s <="111111001010"; -- Argumento 1173 Funcion 0.97399296
  when "010010010110"=> s <="111111001010"; -- Argumento 1174 Funcion 0.97364425
  when "010010010111"=> s <="111111001001"; -- Argumento 1175 Funcion 0.97329325
  when "010010011000"=> s <="111111001000"; -- Argumento 1176 Funcion 0.97293995
  when "010010011001"=> s <="111111000111"; -- Argumento 1177 Funcion 0.97258437
  when "010010011010"=> s <="111111000111"; -- Argumento 1178 Funcion 0.97222650
  when "010010011011"=> s <="111111000110"; -- Argumento 1179 Funcion 0.97186634
  when "010010011100"=> s <="111111000101"; -- Argumento 1180 Funcion 0.97150389
  when "010010011101"=> s <="111111000100"; -- Argumento 1181 Funcion 0.97113916
  when "010010011110"=> s <="111111000100"; -- Argumento 1182 Funcion 0.97077214
  when "010010011111"=> s <="111111000011"; -- Argumento 1183 Funcion 0.97040284
  when "010010100000"=> s <="111111000010"; -- Argumento 1184 Funcion 0.97003125
  when "010010100001"=> s <="111111000001"; -- Argumento 1185 Funcion 0.96965739
  when "010010100010"=> s <="111111000001"; -- Argumento 1186 Funcion 0.96928124
  when "010010100011"=> s <="111111000000"; -- Argumento 1187 Funcion 0.96890280
  when "010010100100"=> s <="111110111111"; -- Argumento 1188 Funcion 0.96852209
  when "010010100101"=> s <="111110111110"; -- Argumento 1189 Funcion 0.96813910
  when "010010100110"=> s <="111110111101"; -- Argumento 1190 Funcion 0.96775384
  when "010010100111"=> s <="111110111101"; -- Argumento 1191 Funcion 0.96736629
  when "010010101000"=> s <="111110111100"; -- Argumento 1192 Funcion 0.96697647
  when "010010101001"=> s <="111110111011"; -- Argumento 1193 Funcion 0.96658437
  when "010010101010"=> s <="111110111010"; -- Argumento 1194 Funcion 0.96619000
  when "010010101011"=> s <="111110111001"; -- Argumento 1195 Funcion 0.96579336
  when "010010101100"=> s <="111110111001"; -- Argumento 1196 Funcion 0.96539444
  when "010010101101"=> s <="111110111000"; -- Argumento 1197 Funcion 0.96499325
  when "010010101110"=> s <="111110110111"; -- Argumento 1198 Funcion 0.96458979
  when "010010101111"=> s <="111110110110"; -- Argumento 1199 Funcion 0.96418406
  when "010010110000"=> s <="111110110101"; -- Argumento 1200 Funcion 0.96377607
  when "010010110001"=> s <="111110110100"; -- Argumento 1201 Funcion 0.96336580
  when "010010110010"=> s <="111110110100"; -- Argumento 1202 Funcion 0.96295327
  when "010010110011"=> s <="111110110011"; -- Argumento 1203 Funcion 0.96253847
  when "010010110100"=> s <="111110110010"; -- Argumento 1204 Funcion 0.96212140
  when "010010110101"=> s <="111110110001"; -- Argumento 1205 Funcion 0.96170208
  when "010010110110"=> s <="111110110000"; -- Argumento 1206 Funcion 0.96128049
  when "010010110111"=> s <="111110101111"; -- Argumento 1207 Funcion 0.96085663
  when "010010111000"=> s <="111110101110"; -- Argumento 1208 Funcion 0.96043052
  when "010010111001"=> s <="111110101110"; -- Argumento 1209 Funcion 0.96000215
  when "010010111010"=> s <="111110101101"; -- Argumento 1210 Funcion 0.95957151
  when "010010111011"=> s <="111110101100"; -- Argumento 1211 Funcion 0.95913862
  when "010010111100"=> s <="111110101011"; -- Argumento 1212 Funcion 0.95870347
  when "010010111101"=> s <="111110101010"; -- Argumento 1213 Funcion 0.95826607
  when "010010111110"=> s <="111110101001"; -- Argumento 1214 Funcion 0.95782641
  when "010010111111"=> s <="111110101000"; -- Argumento 1215 Funcion 0.95738450
  when "010011000000"=> s <="111110100111"; -- Argumento 1216 Funcion 0.95694034
  when "010011000001"=> s <="111110100110"; -- Argumento 1217 Funcion 0.95649392
  when "010011000010"=> s <="111110100101"; -- Argumento 1218 Funcion 0.95604525
  when "010011000011"=> s <="111110100101"; -- Argumento 1219 Funcion 0.95559433
  when "010011000100"=> s <="111110100100"; -- Argumento 1220 Funcion 0.95514117
  when "010011000101"=> s <="111110100011"; -- Argumento 1221 Funcion 0.95468575
  when "010011000110"=> s <="111110100010"; -- Argumento 1222 Funcion 0.95422810
  when "010011000111"=> s <="111110100001"; -- Argumento 1223 Funcion 0.95376819
  when "010011001000"=> s <="111110100000"; -- Argumento 1224 Funcion 0.95330604
  when "010011001001"=> s <="111110011111"; -- Argumento 1225 Funcion 0.95284165
  when "010011001010"=> s <="111110011110"; -- Argumento 1226 Funcion 0.95237501
  when "010011001011"=> s <="111110011101"; -- Argumento 1227 Funcion 0.95190614
  when "010011001100"=> s <="111110011100"; -- Argumento 1228 Funcion 0.95143502
  when "010011001101"=> s <="111110011011"; -- Argumento 1229 Funcion 0.95096167
  when "010011001110"=> s <="111110011010"; -- Argumento 1230 Funcion 0.95048607
  when "010011001111"=> s <="111110011001"; -- Argumento 1231 Funcion 0.95000825
  when "010011010000"=> s <="111110011000"; -- Argumento 1232 Funcion 0.94952818
  when "010011010001"=> s <="111110010111"; -- Argumento 1233 Funcion 0.94904588
  when "010011010010"=> s <="111110010110"; -- Argumento 1234 Funcion 0.94856135
  when "010011010011"=> s <="111110010101"; -- Argumento 1235 Funcion 0.94807459
  when "010011010100"=> s <="111110010100"; -- Argumento 1236 Funcion 0.94758559
  when "010011010101"=> s <="111110010011"; -- Argumento 1237 Funcion 0.94709437
  when "010011010110"=> s <="111110010010"; -- Argumento 1238 Funcion 0.94660091
  when "010011010111"=> s <="111110010001"; -- Argumento 1239 Funcion 0.94610523
  when "010011011000"=> s <="111110010000"; -- Argumento 1240 Funcion 0.94560733
  when "010011011001"=> s <="111110001111"; -- Argumento 1241 Funcion 0.94510719
  when "010011011010"=> s <="111110001110"; -- Argumento 1242 Funcion 0.94460484
  when "010011011011"=> s <="111110001101"; -- Argumento 1243 Funcion 0.94410026
  when "010011011100"=> s <="111110001100"; -- Argumento 1244 Funcion 0.94359346
  when "010011011101"=> s <="111110001011"; -- Argumento 1245 Funcion 0.94308444
  when "010011011110"=> s <="111110001010"; -- Argumento 1246 Funcion 0.94257320
  when "010011011111"=> s <="111110001001"; -- Argumento 1247 Funcion 0.94205974
  when "010011100000"=> s <="111110001000"; -- Argumento 1248 Funcion 0.94154407
  when "010011100001"=> s <="111110000111"; -- Argumento 1249 Funcion 0.94102618
  when "010011100010"=> s <="111110000110"; -- Argumento 1250 Funcion 0.94050607
  when "010011100011"=> s <="111110000101"; -- Argumento 1251 Funcion 0.93998375
  when "010011100100"=> s <="111110000100"; -- Argumento 1252 Funcion 0.93945922
  when "010011100101"=> s <="111110000010"; -- Argumento 1253 Funcion 0.93893248
  when "010011100110"=> s <="111110000001"; -- Argumento 1254 Funcion 0.93840353
  when "010011100111"=> s <="111110000000"; -- Argumento 1255 Funcion 0.93787238
  when "010011101000"=> s <="111101111111"; -- Argumento 1256 Funcion 0.93733901
  when "010011101001"=> s <="111101111110"; -- Argumento 1257 Funcion 0.93680344
  when "010011101010"=> s <="111101111101"; -- Argumento 1258 Funcion 0.93626567
  when "010011101011"=> s <="111101111100"; -- Argumento 1259 Funcion 0.93572569
  when "010011101100"=> s <="111101111011"; -- Argumento 1260 Funcion 0.93518351
  when "010011101101"=> s <="111101111010"; -- Argumento 1261 Funcion 0.93463913
  when "010011101110"=> s <="111101111001"; -- Argumento 1262 Funcion 0.93409255
  when "010011101111"=> s <="111101110111"; -- Argumento 1263 Funcion 0.93354377
  when "010011110000"=> s <="111101110110"; -- Argumento 1264 Funcion 0.93299280
  when "010011110001"=> s <="111101110101"; -- Argumento 1265 Funcion 0.93243963
  when "010011110010"=> s <="111101110100"; -- Argumento 1266 Funcion 0.93188427
  when "010011110011"=> s <="111101110011"; -- Argumento 1267 Funcion 0.93132671
  when "010011110100"=> s <="111101110010"; -- Argumento 1268 Funcion 0.93076696
  when "010011110101"=> s <="111101110001"; -- Argumento 1269 Funcion 0.93020502
  when "010011110110"=> s <="111101101111"; -- Argumento 1270 Funcion 0.92964090
  when "010011110111"=> s <="111101101110"; -- Argumento 1271 Funcion 0.92907458
  when "010011111000"=> s <="111101101101"; -- Argumento 1272 Funcion 0.92850608
  when "010011111001"=> s <="111101101100"; -- Argumento 1273 Funcion 0.92793539
  when "010011111010"=> s <="111101101011"; -- Argumento 1274 Funcion 0.92736253
  when "010011111011"=> s <="111101101010"; -- Argumento 1275 Funcion 0.92678747
  when "010011111100"=> s <="111101101000"; -- Argumento 1276 Funcion 0.92621024
  when "010011111101"=> s <="111101100111"; -- Argumento 1277 Funcion 0.92563083
  when "010011111110"=> s <="111101100110"; -- Argumento 1278 Funcion 0.92504924
  when "010011111111"=> s <="111101100101"; -- Argumento 1279 Funcion 0.92446547
  when "010100000000"=> s <="111101100100"; -- Argumento 1280 Funcion 0.92387953
  when "010100000001"=> s <="111101100010"; -- Argumento 1281 Funcion 0.92329142
  when "010100000010"=> s <="111101100001"; -- Argumento 1282 Funcion 0.92270113
  when "010100000011"=> s <="111101100000"; -- Argumento 1283 Funcion 0.92210867
  when "010100000100"=> s <="111101011111"; -- Argumento 1284 Funcion 0.92151404
  when "010100000101"=> s <="111101011110"; -- Argumento 1285 Funcion 0.92091724
  when "010100000110"=> s <="111101011100"; -- Argumento 1286 Funcion 0.92031828
  when "010100000111"=> s <="111101011011"; -- Argumento 1287 Funcion 0.91971715
  when "010100001000"=> s <="111101011010"; -- Argumento 1288 Funcion 0.91911385
  when "010100001001"=> s <="111101011001"; -- Argumento 1289 Funcion 0.91850839
  when "010100001010"=> s <="111101010111"; -- Argumento 1290 Funcion 0.91790078
  when "010100001011"=> s <="111101010110"; -- Argumento 1291 Funcion 0.91729100
  when "010100001100"=> s <="111101010101"; -- Argumento 1292 Funcion 0.91667906
  when "010100001101"=> s <="111101010100"; -- Argumento 1293 Funcion 0.91606497
  when "010100001110"=> s <="111101010010"; -- Argumento 1294 Funcion 0.91544872
  when "010100001111"=> s <="111101010001"; -- Argumento 1295 Funcion 0.91483031
  when "010100010000"=> s <="111101010000"; -- Argumento 1296 Funcion 0.91420976
  when "010100010001"=> s <="111101001111"; -- Argumento 1297 Funcion 0.91358705
  when "010100010010"=> s <="111101001101"; -- Argumento 1298 Funcion 0.91296219
  when "010100010011"=> s <="111101001100"; -- Argumento 1299 Funcion 0.91233518
  when "010100010100"=> s <="111101001011"; -- Argumento 1300 Funcion 0.91170603
  when "010100010101"=> s <="111101001001"; -- Argumento 1301 Funcion 0.91107473
  when "010100010110"=> s <="111101001000"; -- Argumento 1302 Funcion 0.91044129
  when "010100010111"=> s <="111101000111"; -- Argumento 1303 Funcion 0.90980571
  when "010100011000"=> s <="111101000101"; -- Argumento 1304 Funcion 0.90916798
  when "010100011001"=> s <="111101000100"; -- Argumento 1305 Funcion 0.90852812
  when "010100011010"=> s <="111101000011"; -- Argumento 1306 Funcion 0.90788612
  when "010100011011"=> s <="111101000010"; -- Argumento 1307 Funcion 0.90724198
  when "010100011100"=> s <="111101000000"; -- Argumento 1308 Funcion 0.90659570
  when "010100011101"=> s <="111100111111"; -- Argumento 1309 Funcion 0.90594730
  when "010100011110"=> s <="111100111110"; -- Argumento 1310 Funcion 0.90529676
  when "010100011111"=> s <="111100111100"; -- Argumento 1311 Funcion 0.90464409
  when "010100100000"=> s <="111100111011"; -- Argumento 1312 Funcion 0.90398929
  when "010100100001"=> s <="111100111010"; -- Argumento 1313 Funcion 0.90333237
  when "010100100010"=> s <="111100111000"; -- Argumento 1314 Funcion 0.90267332
  when "010100100011"=> s <="111100110111"; -- Argumento 1315 Funcion 0.90201214
  when "010100100100"=> s <="111100110101"; -- Argumento 1316 Funcion 0.90134885
  when "010100100101"=> s <="111100110100"; -- Argumento 1317 Funcion 0.90068343
  when "010100100110"=> s <="111100110011"; -- Argumento 1318 Funcion 0.90001589
  when "010100100111"=> s <="111100110001"; -- Argumento 1319 Funcion 0.89934624
  when "010100101000"=> s <="111100110000"; -- Argumento 1320 Funcion 0.89867447
  when "010100101001"=> s <="111100101111"; -- Argumento 1321 Funcion 0.89800058
  when "010100101010"=> s <="111100101101"; -- Argumento 1322 Funcion 0.89732458
  when "010100101011"=> s <="111100101100"; -- Argumento 1323 Funcion 0.89664647
  when "010100101100"=> s <="111100101010"; -- Argumento 1324 Funcion 0.89596625
  when "010100101101"=> s <="111100101001"; -- Argumento 1325 Funcion 0.89528392
  when "010100101110"=> s <="111100101000"; -- Argumento 1326 Funcion 0.89459949
  when "010100101111"=> s <="111100100110"; -- Argumento 1327 Funcion 0.89391295
  when "010100110000"=> s <="111100100101"; -- Argumento 1328 Funcion 0.89322430
  when "010100110001"=> s <="111100100011"; -- Argumento 1329 Funcion 0.89253356
  when "010100110010"=> s <="111100100010"; -- Argumento 1330 Funcion 0.89184071
  when "010100110011"=> s <="111100100001"; -- Argumento 1331 Funcion 0.89114576
  when "010100110100"=> s <="111100011111"; -- Argumento 1332 Funcion 0.89044872
  when "010100110101"=> s <="111100011110"; -- Argumento 1333 Funcion 0.88974959
  when "010100110110"=> s <="111100011100"; -- Argumento 1334 Funcion 0.88904836
  when "010100110111"=> s <="111100011011"; -- Argumento 1335 Funcion 0.88834503
  when "010100111000"=> s <="111100011001"; -- Argumento 1336 Funcion 0.88763962
  when "010100111001"=> s <="111100011000"; -- Argumento 1337 Funcion 0.88693212
  when "010100111010"=> s <="111100010110"; -- Argumento 1338 Funcion 0.88622253
  when "010100111011"=> s <="111100010101"; -- Argumento 1339 Funcion 0.88551086
  when "010100111100"=> s <="111100010100"; -- Argumento 1340 Funcion 0.88479710
  when "010100111101"=> s <="111100010010"; -- Argumento 1341 Funcion 0.88408126
  when "010100111110"=> s <="111100010001"; -- Argumento 1342 Funcion 0.88336334
  when "010100111111"=> s <="111100001111"; -- Argumento 1343 Funcion 0.88264334
  when "010101000000"=> s <="111100001110"; -- Argumento 1344 Funcion 0.88192126
  when "010101000001"=> s <="111100001100"; -- Argumento 1345 Funcion 0.88119711
  when "010101000010"=> s <="111100001011"; -- Argumento 1346 Funcion 0.88047089
  when "010101000011"=> s <="111100001001"; -- Argumento 1347 Funcion 0.87974259
  when "010101000100"=> s <="111100001000"; -- Argumento 1348 Funcion 0.87901223
  when "010101000101"=> s <="111100000110"; -- Argumento 1349 Funcion 0.87827979
  when "010101000110"=> s <="111100000101"; -- Argumento 1350 Funcion 0.87754529
  when "010101000111"=> s <="111100000011"; -- Argumento 1351 Funcion 0.87680872
  when "010101001000"=> s <="111100000010"; -- Argumento 1352 Funcion 0.87607009
  when "010101001001"=> s <="111100000000"; -- Argumento 1353 Funcion 0.87532940
  when "010101001010"=> s <="111011111111"; -- Argumento 1354 Funcion 0.87458665
  when "010101001011"=> s <="111011111101"; -- Argumento 1355 Funcion 0.87384184
  when "010101001100"=> s <="111011111100"; -- Argumento 1356 Funcion 0.87309498
  when "010101001101"=> s <="111011111010"; -- Argumento 1357 Funcion 0.87234606
  when "010101001110"=> s <="111011111001"; -- Argumento 1358 Funcion 0.87159509
  when "010101001111"=> s <="111011110111"; -- Argumento 1359 Funcion 0.87084206
  when "010101010000"=> s <="111011110101"; -- Argumento 1360 Funcion 0.87008699
  when "010101010001"=> s <="111011110100"; -- Argumento 1361 Funcion 0.86932987
  when "010101010010"=> s <="111011110010"; -- Argumento 1362 Funcion 0.86857071
  when "010101010011"=> s <="111011110001"; -- Argumento 1363 Funcion 0.86780950
  when "010101010100"=> s <="111011101111"; -- Argumento 1364 Funcion 0.86704625
  when "010101010101"=> s <="111011101110"; -- Argumento 1365 Funcion 0.86628095
  when "010101010110"=> s <="111011101100"; -- Argumento 1366 Funcion 0.86551362
  when "010101010111"=> s <="111011101010"; -- Argumento 1367 Funcion 0.86474426
  when "010101011000"=> s <="111011101001"; -- Argumento 1368 Funcion 0.86397286
  when "010101011001"=> s <="111011100111"; -- Argumento 1369 Funcion 0.86319942
  when "010101011010"=> s <="111011100110"; -- Argumento 1370 Funcion 0.86242396
  when "010101011011"=> s <="111011100100"; -- Argumento 1371 Funcion 0.86164646
  when "010101011100"=> s <="111011100011"; -- Argumento 1372 Funcion 0.86086694
  when "010101011101"=> s <="111011100001"; -- Argumento 1373 Funcion 0.86008539
  when "010101011110"=> s <="111011011111"; -- Argumento 1374 Funcion 0.85930182
  when "010101011111"=> s <="111011011110"; -- Argumento 1375 Funcion 0.85851622
  when "010101100000"=> s <="111011011100"; -- Argumento 1376 Funcion 0.85772861
  when "010101100001"=> s <="111011011011"; -- Argumento 1377 Funcion 0.85693898
  when "010101100010"=> s <="111011011001"; -- Argumento 1378 Funcion 0.85614733
  when "010101100011"=> s <="111011010111"; -- Argumento 1379 Funcion 0.85535366
  when "010101100100"=> s <="111011010110"; -- Argumento 1380 Funcion 0.85455799
  when "010101100101"=> s <="111011010100"; -- Argumento 1381 Funcion 0.85376030
  when "010101100110"=> s <="111011010010"; -- Argumento 1382 Funcion 0.85296060
  when "010101100111"=> s <="111011010001"; -- Argumento 1383 Funcion 0.85215890
  when "010101101000"=> s <="111011001111"; -- Argumento 1384 Funcion 0.85135519
  when "010101101001"=> s <="111011001101"; -- Argumento 1385 Funcion 0.85054948
  when "010101101010"=> s <="111011001100"; -- Argumento 1386 Funcion 0.84974177
  when "010101101011"=> s <="111011001010"; -- Argumento 1387 Funcion 0.84893206
  when "010101101100"=> s <="111011001000"; -- Argumento 1388 Funcion 0.84812034
  when "010101101101"=> s <="111011000111"; -- Argumento 1389 Funcion 0.84730664
  when "010101101110"=> s <="111011000101"; -- Argumento 1390 Funcion 0.84649094
  when "010101101111"=> s <="111011000011"; -- Argumento 1391 Funcion 0.84567325
  when "010101110000"=> s <="111011000010"; -- Argumento 1392 Funcion 0.84485357
  when "010101110001"=> s <="111011000000"; -- Argumento 1393 Funcion 0.84403190
  when "010101110010"=> s <="111010111110"; -- Argumento 1394 Funcion 0.84320824
  when "010101110011"=> s <="111010111101"; -- Argumento 1395 Funcion 0.84238260
  when "010101110100"=> s <="111010111011"; -- Argumento 1396 Funcion 0.84155498
  when "010101110101"=> s <="111010111001"; -- Argumento 1397 Funcion 0.84072537
  when "010101110110"=> s <="111010111000"; -- Argumento 1398 Funcion 0.83989379
  when "010101110111"=> s <="111010110110"; -- Argumento 1399 Funcion 0.83906024
  when "010101111000"=> s <="111010110100"; -- Argumento 1400 Funcion 0.83822471
  when "010101111001"=> s <="111010110010"; -- Argumento 1401 Funcion 0.83738720
  when "010101111010"=> s <="111010110001"; -- Argumento 1402 Funcion 0.83654773
  when "010101111011"=> s <="111010101111"; -- Argumento 1403 Funcion 0.83570628
  when "010101111100"=> s <="111010101101"; -- Argumento 1404 Funcion 0.83486287
  when "010101111101"=> s <="111010101100"; -- Argumento 1405 Funcion 0.83401750
  when "010101111110"=> s <="111010101010"; -- Argumento 1406 Funcion 0.83317016
  when "010101111111"=> s <="111010101000"; -- Argumento 1407 Funcion 0.83232087
  when "010110000000"=> s <="111010100110"; -- Argumento 1408 Funcion 0.83146961
  when "010110000001"=> s <="111010100101"; -- Argumento 1409 Funcion 0.83061640
  when "010110000010"=> s <="111010100011"; -- Argumento 1410 Funcion 0.82976123
  when "010110000011"=> s <="111010100001"; -- Argumento 1411 Funcion 0.82890411
  when "010110000100"=> s <="111010011111"; -- Argumento 1412 Funcion 0.82804505
  when "010110000101"=> s <="111010011110"; -- Argumento 1413 Funcion 0.82718403
  when "010110000110"=> s <="111010011100"; -- Argumento 1414 Funcion 0.82632106
  when "010110000111"=> s <="111010011010"; -- Argumento 1415 Funcion 0.82545615
  when "010110001000"=> s <="111010011000"; -- Argumento 1416 Funcion 0.82458930
  when "010110001001"=> s <="111010010110"; -- Argumento 1417 Funcion 0.82372051
  when "010110001010"=> s <="111010010101"; -- Argumento 1418 Funcion 0.82284978
  when "010110001011"=> s <="111010010011"; -- Argumento 1419 Funcion 0.82197712
  when "010110001100"=> s <="111010010001"; -- Argumento 1420 Funcion 0.82110251
  when "010110001101"=> s <="111010001111"; -- Argumento 1421 Funcion 0.82022598
  when "010110001110"=> s <="111010001110"; -- Argumento 1422 Funcion 0.81934752
  when "010110001111"=> s <="111010001100"; -- Argumento 1423 Funcion 0.81846713
  when "010110010000"=> s <="111010001010"; -- Argumento 1424 Funcion 0.81758481
  when "010110010001"=> s <="111010001000"; -- Argumento 1425 Funcion 0.81670057
  when "010110010010"=> s <="111010000110"; -- Argumento 1426 Funcion 0.81581441
  when "010110010011"=> s <="111010000100"; -- Argumento 1427 Funcion 0.81492633
  when "010110010100"=> s <="111010000011"; -- Argumento 1428 Funcion 0.81403633
  when "010110010101"=> s <="111010000001"; -- Argumento 1429 Funcion 0.81314441
  when "010110010110"=> s <="111001111111"; -- Argumento 1430 Funcion 0.81225059
  when "010110010111"=> s <="111001111101"; -- Argumento 1431 Funcion 0.81135485
  when "010110011000"=> s <="111001111011"; -- Argumento 1432 Funcion 0.81045720
  when "010110011001"=> s <="111001111001"; -- Argumento 1433 Funcion 0.80955764
  when "010110011010"=> s <="111001111000"; -- Argumento 1434 Funcion 0.80865618
  when "010110011011"=> s <="111001110110"; -- Argumento 1435 Funcion 0.80775282
  when "010110011100"=> s <="111001110100"; -- Argumento 1436 Funcion 0.80684755
  when "010110011101"=> s <="111001110010"; -- Argumento 1437 Funcion 0.80594039
  when "010110011110"=> s <="111001110000"; -- Argumento 1438 Funcion 0.80503133
  when "010110011111"=> s <="111001101110"; -- Argumento 1439 Funcion 0.80412038
  when "010110100000"=> s <="111001101100"; -- Argumento 1440 Funcion 0.80320753
  when "010110100001"=> s <="111001101011"; -- Argumento 1441 Funcion 0.80229280
  when "010110100010"=> s <="111001101001"; -- Argumento 1442 Funcion 0.80137617
  when "010110100011"=> s <="111001100111"; -- Argumento 1443 Funcion 0.80045766
  when "010110100100"=> s <="111001100101"; -- Argumento 1444 Funcion 0.79953727
  when "010110100101"=> s <="111001100011"; -- Argumento 1445 Funcion 0.79861499
  when "010110100110"=> s <="111001100001"; -- Argumento 1446 Funcion 0.79769084
  when "010110100111"=> s <="111001011111"; -- Argumento 1447 Funcion 0.79676481
  when "010110101000"=> s <="111001011101"; -- Argumento 1448 Funcion 0.79583690
  when "010110101001"=> s <="111001011011"; -- Argumento 1449 Funcion 0.79490713
  when "010110101010"=> s <="111001011010"; -- Argumento 1450 Funcion 0.79397548
  when "010110101011"=> s <="111001011000"; -- Argumento 1451 Funcion 0.79304196
  when "010110101100"=> s <="111001010110"; -- Argumento 1452 Funcion 0.79210658
  when "010110101101"=> s <="111001010100"; -- Argumento 1453 Funcion 0.79116933
  when "010110101110"=> s <="111001010010"; -- Argumento 1454 Funcion 0.79023022
  when "010110101111"=> s <="111001010000"; -- Argumento 1455 Funcion 0.78928925
  when "010110110000"=> s <="111001001110"; -- Argumento 1456 Funcion 0.78834643
  when "010110110001"=> s <="111001001100"; -- Argumento 1457 Funcion 0.78740175
  when "010110110010"=> s <="111001001010"; -- Argumento 1458 Funcion 0.78645521
  when "010110110011"=> s <="111001001000"; -- Argumento 1459 Funcion 0.78550683
  when "010110110100"=> s <="111001000110"; -- Argumento 1460 Funcion 0.78455660
  when "010110110101"=> s <="111001000100"; -- Argumento 1461 Funcion 0.78360452
  when "010110110110"=> s <="111001000010"; -- Argumento 1462 Funcion 0.78265060
  when "010110110111"=> s <="111001000000"; -- Argumento 1463 Funcion 0.78169483
  when "010110111000"=> s <="111000111110"; -- Argumento 1464 Funcion 0.78073723
  when "010110111001"=> s <="111000111100"; -- Argumento 1465 Funcion 0.77977779
  when "010110111010"=> s <="111000111011"; -- Argumento 1466 Funcion 0.77881651
  when "010110111011"=> s <="111000111001"; -- Argumento 1467 Funcion 0.77785340
  when "010110111100"=> s <="111000110111"; -- Argumento 1468 Funcion 0.77688847
  when "010110111101"=> s <="111000110101"; -- Argumento 1469 Funcion 0.77592170
  when "010110111110"=> s <="111000110011"; -- Argumento 1470 Funcion 0.77495311
  when "010110111111"=> s <="111000110001"; -- Argumento 1471 Funcion 0.77398269
  when "010111000000"=> s <="111000101111"; -- Argumento 1472 Funcion 0.77301045
  when "010111000001"=> s <="111000101101"; -- Argumento 1473 Funcion 0.77203640
  when "010111000010"=> s <="111000101011"; -- Argumento 1474 Funcion 0.77106052
  when "010111000011"=> s <="111000101001"; -- Argumento 1475 Funcion 0.77008284
  when "010111000100"=> s <="111000100111"; -- Argumento 1476 Funcion 0.76910334
  when "010111000101"=> s <="111000100101"; -- Argumento 1477 Funcion 0.76812203
  when "010111000110"=> s <="111000100011"; -- Argumento 1478 Funcion 0.76713891
  when "010111000111"=> s <="111000100001"; -- Argumento 1479 Funcion 0.76615399
  when "010111001000"=> s <="111000011111"; -- Argumento 1480 Funcion 0.76516727
  when "010111001001"=> s <="111000011101"; -- Argumento 1481 Funcion 0.76417874
  when "010111001010"=> s <="111000011011"; -- Argumento 1482 Funcion 0.76318842
  when "010111001011"=> s <="111000011000"; -- Argumento 1483 Funcion 0.76219630
  when "010111001100"=> s <="111000010110"; -- Argumento 1484 Funcion 0.76120239
  when "010111001101"=> s <="111000010100"; -- Argumento 1485 Funcion 0.76020668
  when "010111001110"=> s <="111000010010"; -- Argumento 1486 Funcion 0.75920919
  when "010111001111"=> s <="111000010000"; -- Argumento 1487 Funcion 0.75820991
  when "010111010000"=> s <="111000001110"; -- Argumento 1488 Funcion 0.75720885
  when "010111010001"=> s <="111000001100"; -- Argumento 1489 Funcion 0.75620600
  when "010111010010"=> s <="111000001010"; -- Argumento 1490 Funcion 0.75520138
  when "010111010011"=> s <="111000001000"; -- Argumento 1491 Funcion 0.75419498
  when "010111010100"=> s <="111000000110"; -- Argumento 1492 Funcion 0.75318680
  when "010111010101"=> s <="111000000100"; -- Argumento 1493 Funcion 0.75217685
  when "010111010110"=> s <="111000000010"; -- Argumento 1494 Funcion 0.75116513
  when "010111010111"=> s <="111000000000"; -- Argumento 1495 Funcion 0.75015165
  when "010111011000"=> s <="110111111110"; -- Argumento 1496 Funcion 0.74913639
  when "010111011001"=> s <="110111111100"; -- Argumento 1497 Funcion 0.74811938
  when "010111011010"=> s <="110111111010"; -- Argumento 1498 Funcion 0.74710061
  when "010111011011"=> s <="110111110111"; -- Argumento 1499 Funcion 0.74608007
  when "010111011100"=> s <="110111110101"; -- Argumento 1500 Funcion 0.74505779
  when "010111011101"=> s <="110111110011"; -- Argumento 1501 Funcion 0.74403374
  when "010111011110"=> s <="110111110001"; -- Argumento 1502 Funcion 0.74300795
  when "010111011111"=> s <="110111101111"; -- Argumento 1503 Funcion 0.74198041
  when "010111100000"=> s <="110111101101"; -- Argumento 1504 Funcion 0.74095113
  when "010111100001"=> s <="110111101011"; -- Argumento 1505 Funcion 0.73992010
  when "010111100010"=> s <="110111101001"; -- Argumento 1506 Funcion 0.73888732
  when "010111100011"=> s <="110111100111"; -- Argumento 1507 Funcion 0.73785281
  when "010111100100"=> s <="110111100101"; -- Argumento 1508 Funcion 0.73681657
  when "010111100101"=> s <="110111100010"; -- Argumento 1509 Funcion 0.73577859
  when "010111100110"=> s <="110111100000"; -- Argumento 1510 Funcion 0.73473888
  when "010111100111"=> s <="110111011110"; -- Argumento 1511 Funcion 0.73369744
  when "010111101000"=> s <="110111011100"; -- Argumento 1512 Funcion 0.73265427
  when "010111101001"=> s <="110111011010"; -- Argumento 1513 Funcion 0.73160938
  when "010111101010"=> s <="110111011000"; -- Argumento 1514 Funcion 0.73056277
  when "010111101011"=> s <="110111010110"; -- Argumento 1515 Funcion 0.72951444
  when "010111101100"=> s <="110111010011"; -- Argumento 1516 Funcion 0.72846439
  when "010111101101"=> s <="110111010001"; -- Argumento 1517 Funcion 0.72741263
  when "010111101110"=> s <="110111001111"; -- Argumento 1518 Funcion 0.72635916
  when "010111101111"=> s <="110111001101"; -- Argumento 1519 Funcion 0.72530397
  when "010111110000"=> s <="110111001011"; -- Argumento 1520 Funcion 0.72424708
  when "010111110001"=> s <="110111001001"; -- Argumento 1521 Funcion 0.72318849
  when "010111110010"=> s <="110111000110"; -- Argumento 1522 Funcion 0.72212819
  when "010111110011"=> s <="110111000100"; -- Argumento 1523 Funcion 0.72106620
  when "010111110100"=> s <="110111000010"; -- Argumento 1524 Funcion 0.72000251
  when "010111110101"=> s <="110111000000"; -- Argumento 1525 Funcion 0.71893712
  when "010111110110"=> s <="110110111110"; -- Argumento 1526 Funcion 0.71787005
  when "010111110111"=> s <="110110111100"; -- Argumento 1527 Funcion 0.71680128
  when "010111111000"=> s <="110110111001"; -- Argumento 1528 Funcion 0.71573083
  when "010111111001"=> s <="110110110111"; -- Argumento 1529 Funcion 0.71465869
  when "010111111010"=> s <="110110110101"; -- Argumento 1530 Funcion 0.71358487
  when "010111111011"=> s <="110110110011"; -- Argumento 1531 Funcion 0.71250937
  when "010111111100"=> s <="110110110001"; -- Argumento 1532 Funcion 0.71143220
  when "010111111101"=> s <="110110101110"; -- Argumento 1533 Funcion 0.71035335
  when "010111111110"=> s <="110110101100"; -- Argumento 1534 Funcion 0.70927283
  when "010111111111"=> s <="110110101010"; -- Argumento 1535 Funcion 0.70819064
  when "011000000000"=> s <="110110101000"; -- Argumento 1536 Funcion 0.70710678
  when "011000000001"=> s <="110110100101"; -- Argumento 1537 Funcion 0.70602126
  when "011000000010"=> s <="110110100011"; -- Argumento 1538 Funcion 0.70493408
  when "011000000011"=> s <="110110100001"; -- Argumento 1539 Funcion 0.70384524
  when "011000000100"=> s <="110110011111"; -- Argumento 1540 Funcion 0.70275474
  when "011000000101"=> s <="110110011101"; -- Argumento 1541 Funcion 0.70166259
  when "011000000110"=> s <="110110011010"; -- Argumento 1542 Funcion 0.70056879
  when "011000000111"=> s <="110110011000"; -- Argumento 1543 Funcion 0.69947334
  when "011000001000"=> s <="110110010110"; -- Argumento 1544 Funcion 0.69837625
  when "011000001001"=> s <="110110010100"; -- Argumento 1545 Funcion 0.69727751
  when "011000001010"=> s <="110110010001"; -- Argumento 1546 Funcion 0.69617713
  when "011000001011"=> s <="110110001111"; -- Argumento 1547 Funcion 0.69507511
  when "011000001100"=> s <="110110001101"; -- Argumento 1548 Funcion 0.69397146
  when "011000001101"=> s <="110110001010"; -- Argumento 1549 Funcion 0.69286617
  when "011000001110"=> s <="110110001000"; -- Argumento 1550 Funcion 0.69175926
  when "011000001111"=> s <="110110000110"; -- Argumento 1551 Funcion 0.69065071
  when "011000010000"=> s <="110110000100"; -- Argumento 1552 Funcion 0.68954054
  when "011000010001"=> s <="110110000001"; -- Argumento 1553 Funcion 0.68842875
  when "011000010010"=> s <="110101111111"; -- Argumento 1554 Funcion 0.68731534
  when "011000010011"=> s <="110101111101"; -- Argumento 1555 Funcion 0.68620031
  when "011000010100"=> s <="110101111011"; -- Argumento 1556 Funcion 0.68508367
  when "011000010101"=> s <="110101111000"; -- Argumento 1557 Funcion 0.68396541
  when "011000010110"=> s <="110101110110"; -- Argumento 1558 Funcion 0.68284555
  when "011000010111"=> s <="110101110100"; -- Argumento 1559 Funcion 0.68172407
  when "011000011000"=> s <="110101110001"; -- Argumento 1560 Funcion 0.68060100
  when "011000011001"=> s <="110101101111"; -- Argumento 1561 Funcion 0.67947632
  when "011000011010"=> s <="110101101101"; -- Argumento 1562 Funcion 0.67835004
  when "011000011011"=> s <="110101101010"; -- Argumento 1563 Funcion 0.67722217
  when "011000011100"=> s <="110101101000"; -- Argumento 1564 Funcion 0.67609270
  when "011000011101"=> s <="110101100110"; -- Argumento 1565 Funcion 0.67496165
  when "011000011110"=> s <="110101100100"; -- Argumento 1566 Funcion 0.67382900
  when "011000011111"=> s <="110101100001"; -- Argumento 1567 Funcion 0.67269477
  when "011000100000"=> s <="110101011111"; -- Argumento 1568 Funcion 0.67155895
  when "011000100001"=> s <="110101011101"; -- Argumento 1569 Funcion 0.67042156
  when "011000100010"=> s <="110101011010"; -- Argumento 1570 Funcion 0.66928259
  when "011000100011"=> s <="110101011000"; -- Argumento 1571 Funcion 0.66814204
  when "011000100100"=> s <="110101010110"; -- Argumento 1572 Funcion 0.66699992
  when "011000100101"=> s <="110101010011"; -- Argumento 1573 Funcion 0.66585623
  when "011000100110"=> s <="110101010001"; -- Argumento 1574 Funcion 0.66471098
  when "011000100111"=> s <="110101001110"; -- Argumento 1575 Funcion 0.66356416
  when "011000101000"=> s <="110101001100"; -- Argumento 1576 Funcion 0.66241578
  when "011000101001"=> s <="110101001010"; -- Argumento 1577 Funcion 0.66126584
  when "011000101010"=> s <="110101000111"; -- Argumento 1578 Funcion 0.66011434
  when "011000101011"=> s <="110101000101"; -- Argumento 1579 Funcion 0.65896129
  when "011000101100"=> s <="110101000011"; -- Argumento 1580 Funcion 0.65780669
  when "011000101101"=> s <="110101000000"; -- Argumento 1581 Funcion 0.65665055
  when "011000101110"=> s <="110100111110"; -- Argumento 1582 Funcion 0.65549285
  when "011000101111"=> s <="110100111100"; -- Argumento 1583 Funcion 0.65433362
  when "011000110000"=> s <="110100111001"; -- Argumento 1584 Funcion 0.65317284
  when "011000110001"=> s <="110100110111"; -- Argumento 1585 Funcion 0.65201053
  when "011000110010"=> s <="110100110100"; -- Argumento 1586 Funcion 0.65084668
  when "011000110011"=> s <="110100110010"; -- Argumento 1587 Funcion 0.64968131
  when "011000110100"=> s <="110100110000"; -- Argumento 1588 Funcion 0.64851440
  when "011000110101"=> s <="110100101101"; -- Argumento 1589 Funcion 0.64734597
  when "011000110110"=> s <="110100101011"; -- Argumento 1590 Funcion 0.64617601
  when "011000110111"=> s <="110100101000"; -- Argumento 1591 Funcion 0.64500454
  when "011000111000"=> s <="110100100110"; -- Argumento 1592 Funcion 0.64383154
  when "011000111001"=> s <="110100100100"; -- Argumento 1593 Funcion 0.64265703
  when "011000111010"=> s <="110100100001"; -- Argumento 1594 Funcion 0.64148101
  when "011000111011"=> s <="110100011111"; -- Argumento 1595 Funcion 0.64030348
  when "011000111100"=> s <="110100011100"; -- Argumento 1596 Funcion 0.63912444
  when "011000111101"=> s <="110100011010"; -- Argumento 1597 Funcion 0.63794390
  when "011000111110"=> s <="110100011000"; -- Argumento 1598 Funcion 0.63676186
  when "011000111111"=> s <="110100010101"; -- Argumento 1599 Funcion 0.63557832
  when "011001000000"=> s <="110100010011"; -- Argumento 1600 Funcion 0.63439328
  when "011001000001"=> s <="110100010000"; -- Argumento 1601 Funcion 0.63320676
  when "011001000010"=> s <="110100001110"; -- Argumento 1602 Funcion 0.63201874
  when "011001000011"=> s <="110100001011"; -- Argumento 1603 Funcion 0.63082923
  when "011001000100"=> s <="110100001001"; -- Argumento 1604 Funcion 0.62963824
  when "011001000101"=> s <="110100000111"; -- Argumento 1605 Funcion 0.62844577
  when "011001000110"=> s <="110100000100"; -- Argumento 1606 Funcion 0.62725182
  when "011001000111"=> s <="110100000010"; -- Argumento 1607 Funcion 0.62605639
  when "011001001000"=> s <="110011111111"; -- Argumento 1608 Funcion 0.62485949
  when "011001001001"=> s <="110011111101"; -- Argumento 1609 Funcion 0.62366112
  when "011001001010"=> s <="110011111010"; -- Argumento 1610 Funcion 0.62246128
  when "011001001011"=> s <="110011111000"; -- Argumento 1611 Funcion 0.62125998
  when "011001001100"=> s <="110011110101"; -- Argumento 1612 Funcion 0.62005721
  when "011001001101"=> s <="110011110011"; -- Argumento 1613 Funcion 0.61885299
  when "011001001110"=> s <="110011110000"; -- Argumento 1614 Funcion 0.61764731
  when "011001001111"=> s <="110011101110"; -- Argumento 1615 Funcion 0.61644017
  when "011001010000"=> s <="110011101011"; -- Argumento 1616 Funcion 0.61523159
  when "011001010001"=> s <="110011101001"; -- Argumento 1617 Funcion 0.61402156
  when "011001010010"=> s <="110011100111"; -- Argumento 1618 Funcion 0.61281008
  when "011001010011"=> s <="110011100100"; -- Argumento 1619 Funcion 0.61159716
  when "011001010100"=> s <="110011100010"; -- Argumento 1620 Funcion 0.61038281
  when "011001010101"=> s <="110011011111"; -- Argumento 1621 Funcion 0.60916701
  when "011001010110"=> s <="110011011101"; -- Argumento 1622 Funcion 0.60794978
  when "011001010111"=> s <="110011011010"; -- Argumento 1623 Funcion 0.60673113
  when "011001011000"=> s <="110011011000"; -- Argumento 1624 Funcion 0.60551104
  when "011001011001"=> s <="110011010101"; -- Argumento 1625 Funcion 0.60428953
  when "011001011010"=> s <="110011010011"; -- Argumento 1626 Funcion 0.60306660
  when "011001011011"=> s <="110011010000"; -- Argumento 1627 Funcion 0.60184225
  when "011001011100"=> s <="110011001110"; -- Argumento 1628 Funcion 0.60061648
  when "011001011101"=> s <="110011001011"; -- Argumento 1629 Funcion 0.59938930
  when "011001011110"=> s <="110011001001"; -- Argumento 1630 Funcion 0.59816071
  when "011001011111"=> s <="110011000110"; -- Argumento 1631 Funcion 0.59693071
  when "011001100000"=> s <="110011000011"; -- Argumento 1632 Funcion 0.59569930
  when "011001100001"=> s <="110011000001"; -- Argumento 1633 Funcion 0.59446650
  when "011001100010"=> s <="110010111110"; -- Argumento 1634 Funcion 0.59323230
  when "011001100011"=> s <="110010111100"; -- Argumento 1635 Funcion 0.59199669
  when "011001100100"=> s <="110010111001"; -- Argumento 1636 Funcion 0.59075970
  when "011001100101"=> s <="110010110111"; -- Argumento 1637 Funcion 0.58952132
  when "011001100110"=> s <="110010110100"; -- Argumento 1638 Funcion 0.58828155
  when "011001100111"=> s <="110010110010"; -- Argumento 1639 Funcion 0.58704039
  when "011001101000"=> s <="110010101111"; -- Argumento 1640 Funcion 0.58579786
  when "011001101001"=> s <="110010101101"; -- Argumento 1641 Funcion 0.58455394
  when "011001101010"=> s <="110010101010"; -- Argumento 1642 Funcion 0.58330865
  when "011001101011"=> s <="110010101000"; -- Argumento 1643 Funcion 0.58206199
  when "011001101100"=> s <="110010100101"; -- Argumento 1644 Funcion 0.58081396
  when "011001101101"=> s <="110010100010"; -- Argumento 1645 Funcion 0.57956456
  when "011001101110"=> s <="110010100000"; -- Argumento 1646 Funcion 0.57831380
  when "011001101111"=> s <="110010011101"; -- Argumento 1647 Funcion 0.57706167
  when "011001110000"=> s <="110010011011"; -- Argumento 1648 Funcion 0.57580819
  when "011001110001"=> s <="110010011000"; -- Argumento 1649 Funcion 0.57455336
  when "011001110010"=> s <="110010010110"; -- Argumento 1650 Funcion 0.57329717
  when "011001110011"=> s <="110010010011"; -- Argumento 1651 Funcion 0.57203963
  when "011001110100"=> s <="110010010000"; -- Argumento 1652 Funcion 0.57078075
  when "011001110101"=> s <="110010001110"; -- Argumento 1653 Funcion 0.56952052
  when "011001110110"=> s <="110010001011"; -- Argumento 1654 Funcion 0.56825895
  when "011001110111"=> s <="110010001001"; -- Argumento 1655 Funcion 0.56699605
  when "011001111000"=> s <="110010000110"; -- Argumento 1656 Funcion 0.56573181
  when "011001111001"=> s <="110010000100"; -- Argumento 1657 Funcion 0.56446624
  when "011001111010"=> s <="110010000001"; -- Argumento 1658 Funcion 0.56319934
  when "011001111011"=> s <="110001111110"; -- Argumento 1659 Funcion 0.56193112
  when "011001111100"=> s <="110001111100"; -- Argumento 1660 Funcion 0.56066158
  when "011001111101"=> s <="110001111001"; -- Argumento 1661 Funcion 0.55939071
  when "011001111110"=> s <="110001110111"; -- Argumento 1662 Funcion 0.55811853
  when "011001111111"=> s <="110001110100"; -- Argumento 1663 Funcion 0.55684504
  when "011010000000"=> s <="110001110001"; -- Argumento 1664 Funcion 0.55557023
  when "011010000001"=> s <="110001101111"; -- Argumento 1665 Funcion 0.55429412
  when "011010000010"=> s <="110001101100"; -- Argumento 1666 Funcion 0.55301671
  when "011010000011"=> s <="110001101001"; -- Argumento 1667 Funcion 0.55173799
  when "011010000100"=> s <="110001100111"; -- Argumento 1668 Funcion 0.55045797
  when "011010000101"=> s <="110001100100"; -- Argumento 1669 Funcion 0.54917666
  when "011010000110"=> s <="110001100010"; -- Argumento 1670 Funcion 0.54789406
  when "011010000111"=> s <="110001011111"; -- Argumento 1671 Funcion 0.54661017
  when "011010001000"=> s <="110001011100"; -- Argumento 1672 Funcion 0.54532499
  when "011010001001"=> s <="110001011010"; -- Argumento 1673 Funcion 0.54403853
  when "011010001010"=> s <="110001010111"; -- Argumento 1674 Funcion 0.54275078
  when "011010001011"=> s <="110001010100"; -- Argumento 1675 Funcion 0.54146177
  when "011010001100"=> s <="110001010010"; -- Argumento 1676 Funcion 0.54017147
  when "011010001101"=> s <="110001001111"; -- Argumento 1677 Funcion 0.53887991
  when "011010001110"=> s <="110001001100"; -- Argumento 1678 Funcion 0.53758708
  when "011010001111"=> s <="110001001010"; -- Argumento 1679 Funcion 0.53629298
  when "011010010000"=> s <="110001000111"; -- Argumento 1680 Funcion 0.53499762
  when "011010010001"=> s <="110001000101"; -- Argumento 1681 Funcion 0.53370100
  when "011010010010"=> s <="110001000010"; -- Argumento 1682 Funcion 0.53240313
  when "011010010011"=> s <="110000111111"; -- Argumento 1683 Funcion 0.53110400
  when "011010010100"=> s <="110000111101"; -- Argumento 1684 Funcion 0.52980362
  when "011010010101"=> s <="110000111010"; -- Argumento 1685 Funcion 0.52850200
  when "011010010110"=> s <="110000110111"; -- Argumento 1686 Funcion 0.52719913
  when "011010010111"=> s <="110000110101"; -- Argumento 1687 Funcion 0.52589503
  when "011010011000"=> s <="110000110010"; -- Argumento 1688 Funcion 0.52458968
  when "011010011001"=> s <="110000101111"; -- Argumento 1689 Funcion 0.52328310
  when "011010011010"=> s <="110000101101"; -- Argumento 1690 Funcion 0.52197529
  when "011010011011"=> s <="110000101010"; -- Argumento 1691 Funcion 0.52066625
  when "011010011100"=> s <="110000100111"; -- Argumento 1692 Funcion 0.51935599
  when "011010011101"=> s <="110000100100"; -- Argumento 1693 Funcion 0.51804450
  when "011010011110"=> s <="110000100010"; -- Argumento 1694 Funcion 0.51673180
  when "011010011111"=> s <="110000011111"; -- Argumento 1695 Funcion 0.51541788
  when "011010100000"=> s <="110000011100"; -- Argumento 1696 Funcion 0.51410274
  when "011010100001"=> s <="110000011010"; -- Argumento 1697 Funcion 0.51278640
  when "011010100010"=> s <="110000010111"; -- Argumento 1698 Funcion 0.51146885
  when "011010100011"=> s <="110000010100"; -- Argumento 1699 Funcion 0.51015010
  when "011010100100"=> s <="110000010010"; -- Argumento 1700 Funcion 0.50883014
  when "011010100101"=> s <="110000001111"; -- Argumento 1701 Funcion 0.50750899
  when "011010100110"=> s <="110000001100"; -- Argumento 1702 Funcion 0.50618665
  when "011010100111"=> s <="110000001001"; -- Argumento 1703 Funcion 0.50486311
  when "011010101000"=> s <="110000000111"; -- Argumento 1704 Funcion 0.50353838
  when "011010101001"=> s <="110000000100"; -- Argumento 1705 Funcion 0.50221247
  when "011010101010"=> s <="110000000001"; -- Argumento 1706 Funcion 0.50088538
  when "011010101011"=> s <="101111111111"; -- Argumento 1707 Funcion 0.49955711
  when "011010101100"=> s <="101111111100"; -- Argumento 1708 Funcion 0.49822767
  when "011010101101"=> s <="101111111001"; -- Argumento 1709 Funcion 0.49689705
  when "011010101110"=> s <="101111110110"; -- Argumento 1710 Funcion 0.49556526
  when "011010101111"=> s <="101111110100"; -- Argumento 1711 Funcion 0.49423231
  when "011010110000"=> s <="101111110001"; -- Argumento 1712 Funcion 0.49289819
  when "011010110001"=> s <="101111101110"; -- Argumento 1713 Funcion 0.49156292
  when "011010110010"=> s <="101111101011"; -- Argumento 1714 Funcion 0.49022648
  when "011010110011"=> s <="101111101001"; -- Argumento 1715 Funcion 0.48888890
  when "011010110100"=> s <="101111100110"; -- Argumento 1716 Funcion 0.48755016
  when "011010110101"=> s <="101111100011"; -- Argumento 1717 Funcion 0.48621028
  when "011010110110"=> s <="101111100001"; -- Argumento 1718 Funcion 0.48486925
  when "011010110111"=> s <="101111011110"; -- Argumento 1719 Funcion 0.48352708
  when "011010111000"=> s <="101111011011"; -- Argumento 1720 Funcion 0.48218377
  when "011010111001"=> s <="101111011000"; -- Argumento 1721 Funcion 0.48083933
  when "011010111010"=> s <="101111010110"; -- Argumento 1722 Funcion 0.47949376
  when "011010111011"=> s <="101111010011"; -- Argumento 1723 Funcion 0.47814706
  when "011010111100"=> s <="101111010000"; -- Argumento 1724 Funcion 0.47679923
  when "011010111101"=> s <="101111001101"; -- Argumento 1725 Funcion 0.47545028
  when "011010111110"=> s <="101111001010"; -- Argumento 1726 Funcion 0.47410021
  when "011010111111"=> s <="101111001000"; -- Argumento 1727 Funcion 0.47274903
  when "011011000000"=> s <="101111000101"; -- Argumento 1728 Funcion 0.47139674
  when "011011000001"=> s <="101111000010"; -- Argumento 1729 Funcion 0.47004333
  when "011011000010"=> s <="101110111111"; -- Argumento 1730 Funcion 0.46868882
  when "011011000011"=> s <="101110111101"; -- Argumento 1731 Funcion 0.46733321
  when "011011000100"=> s <="101110111010"; -- Argumento 1732 Funcion 0.46597650
  when "011011000101"=> s <="101110110111"; -- Argumento 1733 Funcion 0.46461869
  when "011011000110"=> s <="101110110100"; -- Argumento 1734 Funcion 0.46325978
  when "011011000111"=> s <="101110110001"; -- Argumento 1735 Funcion 0.46189979
  when "011011001000"=> s <="101110101111"; -- Argumento 1736 Funcion 0.46053871
  when "011011001001"=> s <="101110101100"; -- Argumento 1737 Funcion 0.45917655
  when "011011001010"=> s <="101110101001"; -- Argumento 1738 Funcion 0.45781330
  when "011011001011"=> s <="101110100110"; -- Argumento 1739 Funcion 0.45644898
  when "011011001100"=> s <="101110100100"; -- Argumento 1740 Funcion 0.45508359
  when "011011001101"=> s <="101110100001"; -- Argumento 1741 Funcion 0.45371712
  when "011011001110"=> s <="101110011110"; -- Argumento 1742 Funcion 0.45234959
  when "011011001111"=> s <="101110011011"; -- Argumento 1743 Funcion 0.45098099
  when "011011010000"=> s <="101110011000"; -- Argumento 1744 Funcion 0.44961133
  when "011011010001"=> s <="101110010101"; -- Argumento 1745 Funcion 0.44824061
  when "011011010010"=> s <="101110010011"; -- Argumento 1746 Funcion 0.44686884
  when "011011010011"=> s <="101110010000"; -- Argumento 1747 Funcion 0.44549602
  when "011011010100"=> s <="101110001101"; -- Argumento 1748 Funcion 0.44412214
  when "011011010101"=> s <="101110001010"; -- Argumento 1749 Funcion 0.44274723
  when "011011010110"=> s <="101110000111"; -- Argumento 1750 Funcion 0.44137127
  when "011011010111"=> s <="101110000101"; -- Argumento 1751 Funcion 0.43999427
  when "011011011000"=> s <="101110000010"; -- Argumento 1752 Funcion 0.43861624
  when "011011011001"=> s <="101101111111"; -- Argumento 1753 Funcion 0.43723717
  when "011011011010"=> s <="101101111100"; -- Argumento 1754 Funcion 0.43585708
  when "011011011011"=> s <="101101111001"; -- Argumento 1755 Funcion 0.43447596
  when "011011011100"=> s <="101101110110"; -- Argumento 1756 Funcion 0.43309382
  when "011011011101"=> s <="101101110100"; -- Argumento 1757 Funcion 0.43171066
  when "011011011110"=> s <="101101110001"; -- Argumento 1758 Funcion 0.43032648
  when "011011011111"=> s <="101101101110"; -- Argumento 1759 Funcion 0.42894129
  when "011011100000"=> s <="101101101011"; -- Argumento 1760 Funcion 0.42755509
  when "011011100001"=> s <="101101101000"; -- Argumento 1761 Funcion 0.42616789
  when "011011100010"=> s <="101101100101"; -- Argumento 1762 Funcion 0.42477968
  when "011011100011"=> s <="101101100011"; -- Argumento 1763 Funcion 0.42339047
  when "011011100100"=> s <="101101100000"; -- Argumento 1764 Funcion 0.42200027
  when "011011100101"=> s <="101101011101"; -- Argumento 1765 Funcion 0.42060907
  when "011011100110"=> s <="101101011010"; -- Argumento 1766 Funcion 0.41921689
  when "011011100111"=> s <="101101010111"; -- Argumento 1767 Funcion 0.41782372
  when "011011101000"=> s <="101101010100"; -- Argumento 1768 Funcion 0.41642956
  when "011011101001"=> s <="101101010001"; -- Argumento 1769 Funcion 0.41503442
  when "011011101010"=> s <="101101001111"; -- Argumento 1770 Funcion 0.41363831
  when "011011101011"=> s <="101101001100"; -- Argumento 1771 Funcion 0.41224123
  when "011011101100"=> s <="101101001001"; -- Argumento 1772 Funcion 0.41084317
  when "011011101101"=> s <="101101000110"; -- Argumento 1773 Funcion 0.40944415
  when "011011101110"=> s <="101101000011"; -- Argumento 1774 Funcion 0.40804416
  when "011011101111"=> s <="101101000000"; -- Argumento 1775 Funcion 0.40664322
  when "011011110000"=> s <="101100111101"; -- Argumento 1776 Funcion 0.40524131
  when "011011110001"=> s <="101100111011"; -- Argumento 1777 Funcion 0.40383846
  when "011011110010"=> s <="101100111000"; -- Argumento 1778 Funcion 0.40243465
  when "011011110011"=> s <="101100110101"; -- Argumento 1779 Funcion 0.40102990
  when "011011110100"=> s <="101100110010"; -- Argumento 1780 Funcion 0.39962420
  when "011011110101"=> s <="101100101111"; -- Argumento 1781 Funcion 0.39821756
  when "011011110110"=> s <="101100101100"; -- Argumento 1782 Funcion 0.39680999
  when "011011110111"=> s <="101100101001"; -- Argumento 1783 Funcion 0.39540148
  when "011011111000"=> s <="101100100110"; -- Argumento 1784 Funcion 0.39399204
  when "011011111001"=> s <="101100100100"; -- Argumento 1785 Funcion 0.39258167
  when "011011111010"=> s <="101100100001"; -- Argumento 1786 Funcion 0.39117038
  when "011011111011"=> s <="101100011110"; -- Argumento 1787 Funcion 0.38975817
  when "011011111100"=> s <="101100011011"; -- Argumento 1788 Funcion 0.38834505
  when "011011111101"=> s <="101100011000"; -- Argumento 1789 Funcion 0.38693101
  when "011011111110"=> s <="101100010101"; -- Argumento 1790 Funcion 0.38551605
  when "011011111111"=> s <="101100010010"; -- Argumento 1791 Funcion 0.38410020
  when "011100000000"=> s <="101100001111"; -- Argumento 1792 Funcion 0.38268343
  when "011100000001"=> s <="101100001100"; -- Argumento 1793 Funcion 0.38126577
  when "011100000010"=> s <="101100001001"; -- Argumento 1794 Funcion 0.37984721
  when "011100000011"=> s <="101100000111"; -- Argumento 1795 Funcion 0.37842775
  when "011100000100"=> s <="101100000100"; -- Argumento 1796 Funcion 0.37700741
  when "011100000101"=> s <="101100000001"; -- Argumento 1797 Funcion 0.37558618
  when "011100000110"=> s <="101011111110"; -- Argumento 1798 Funcion 0.37416406
  when "011100000111"=> s <="101011111011"; -- Argumento 1799 Funcion 0.37274107
  when "011100001000"=> s <="101011111000"; -- Argumento 1800 Funcion 0.37131719
  when "011100001001"=> s <="101011110101"; -- Argumento 1801 Funcion 0.36989245
  when "011100001010"=> s <="101011110010"; -- Argumento 1802 Funcion 0.36846683
  when "011100001011"=> s <="101011101111"; -- Argumento 1803 Funcion 0.36704035
  when "011100001100"=> s <="101011101100"; -- Argumento 1804 Funcion 0.36561300
  when "011100001101"=> s <="101011101001"; -- Argumento 1805 Funcion 0.36418479
  when "011100001110"=> s <="101011100110"; -- Argumento 1806 Funcion 0.36275572
  when "011100001111"=> s <="101011100011"; -- Argumento 1807 Funcion 0.36132581
  when "011100010000"=> s <="101011100001"; -- Argumento 1808 Funcion 0.35989504
  when "011100010001"=> s <="101011011110"; -- Argumento 1809 Funcion 0.35846342
  when "011100010010"=> s <="101011011011"; -- Argumento 1810 Funcion 0.35703096
  when "011100010011"=> s <="101011011000"; -- Argumento 1811 Funcion 0.35559766
  when "011100010100"=> s <="101011010101"; -- Argumento 1812 Funcion 0.35416353
  when "011100010101"=> s <="101011010010"; -- Argumento 1813 Funcion 0.35272856
  when "011100010110"=> s <="101011001111"; -- Argumento 1814 Funcion 0.35129276
  when "011100010111"=> s <="101011001100"; -- Argumento 1815 Funcion 0.34985613
  when "011100011000"=> s <="101011001001"; -- Argumento 1816 Funcion 0.34841868
  when "011100011001"=> s <="101011000110"; -- Argumento 1817 Funcion 0.34698041
  when "011100011010"=> s <="101011000011"; -- Argumento 1818 Funcion 0.34554132
  when "011100011011"=> s <="101011000000"; -- Argumento 1819 Funcion 0.34410143
  when "011100011100"=> s <="101010111101"; -- Argumento 1820 Funcion 0.34266072
  when "011100011101"=> s <="101010111010"; -- Argumento 1821 Funcion 0.34121920
  when "011100011110"=> s <="101010110111"; -- Argumento 1822 Funcion 0.33977688
  when "011100011111"=> s <="101010110100"; -- Argumento 1823 Funcion 0.33833377
  when "011100100000"=> s <="101010110001"; -- Argumento 1824 Funcion 0.33688985
  when "011100100001"=> s <="101010101110"; -- Argumento 1825 Funcion 0.33544515
  when "011100100010"=> s <="101010101100"; -- Argumento 1826 Funcion 0.33399965
  when "011100100011"=> s <="101010101001"; -- Argumento 1827 Funcion 0.33255337
  when "011100100100"=> s <="101010100110"; -- Argumento 1828 Funcion 0.33110631
  when "011100100101"=> s <="101010100011"; -- Argumento 1829 Funcion 0.32965846
  when "011100100110"=> s <="101010100000"; -- Argumento 1830 Funcion 0.32820984
  when "011100100111"=> s <="101010011101"; -- Argumento 1831 Funcion 0.32676045
  when "011100101000"=> s <="101010011010"; -- Argumento 1832 Funcion 0.32531029
  when "011100101001"=> s <="101010010111"; -- Argumento 1833 Funcion 0.32385937
  when "011100101010"=> s <="101010010100"; -- Argumento 1834 Funcion 0.32240768
  when "011100101011"=> s <="101010010001"; -- Argumento 1835 Funcion 0.32095523
  when "011100101100"=> s <="101010001110"; -- Argumento 1836 Funcion 0.31950203
  when "011100101101"=> s <="101010001011"; -- Argumento 1837 Funcion 0.31804808
  when "011100101110"=> s <="101010001000"; -- Argumento 1838 Funcion 0.31659338
  when "011100101111"=> s <="101010000101"; -- Argumento 1839 Funcion 0.31513793
  when "011100110000"=> s <="101010000010"; -- Argumento 1840 Funcion 0.31368174
  when "011100110001"=> s <="101001111111"; -- Argumento 1841 Funcion 0.31222481
  when "011100110010"=> s <="101001111100"; -- Argumento 1842 Funcion 0.31076715
  when "011100110011"=> s <="101001111001"; -- Argumento 1843 Funcion 0.30930876
  when "011100110100"=> s <="101001110110"; -- Argumento 1844 Funcion 0.30784964
  when "011100110101"=> s <="101001110011"; -- Argumento 1845 Funcion 0.30638980
  when "011100110110"=> s <="101001110000"; -- Argumento 1846 Funcion 0.30492923
  when "011100110111"=> s <="101001101101"; -- Argumento 1847 Funcion 0.30346795
  when "011100111000"=> s <="101001101010"; -- Argumento 1848 Funcion 0.30200595
  when "011100111001"=> s <="101001100111"; -- Argumento 1849 Funcion 0.30054324
  when "011100111010"=> s <="101001100100"; -- Argumento 1850 Funcion 0.29907983
  when "011100111011"=> s <="101001100001"; -- Argumento 1851 Funcion 0.29761571
  when "011100111100"=> s <="101001011110"; -- Argumento 1852 Funcion 0.29615089
  when "011100111101"=> s <="101001011011"; -- Argumento 1853 Funcion 0.29468537
  when "011100111110"=> s <="101001011000"; -- Argumento 1854 Funcion 0.29321916
  when "011100111111"=> s <="101001010101"; -- Argumento 1855 Funcion 0.29175226
  when "011101000000"=> s <="101001010010"; -- Argumento 1856 Funcion 0.29028468
  when "011101000001"=> s <="101001001111"; -- Argumento 1857 Funcion 0.28881641
  when "011101000010"=> s <="101001001100"; -- Argumento 1858 Funcion 0.28734746
  when "011101000011"=> s <="101001001001"; -- Argumento 1859 Funcion 0.28587783
  when "011101000100"=> s <="101001000110"; -- Argumento 1860 Funcion 0.28440754
  when "011101000101"=> s <="101001000011"; -- Argumento 1861 Funcion 0.28293657
  when "011101000110"=> s <="101001000000"; -- Argumento 1862 Funcion 0.28146494
  when "011101000111"=> s <="101000111101"; -- Argumento 1863 Funcion 0.27999264
  when "011101001000"=> s <="101000111010"; -- Argumento 1864 Funcion 0.27851969
  when "011101001001"=> s <="101000110111"; -- Argumento 1865 Funcion 0.27704608
  when "011101001010"=> s <="101000110100"; -- Argumento 1866 Funcion 0.27557182
  when "011101001011"=> s <="101000110001"; -- Argumento 1867 Funcion 0.27409691
  when "011101001100"=> s <="101000101110"; -- Argumento 1868 Funcion 0.27262136
  when "011101001101"=> s <="101000101011"; -- Argumento 1869 Funcion 0.27114516
  when "011101001110"=> s <="101000101000"; -- Argumento 1870 Funcion 0.26966833
  when "011101001111"=> s <="101000100101"; -- Argumento 1871 Funcion 0.26819086
  when "011101010000"=> s <="101000100010"; -- Argumento 1872 Funcion 0.26671276
  when "011101010001"=> s <="101000011111"; -- Argumento 1873 Funcion 0.26523403
  when "011101010010"=> s <="101000011100"; -- Argumento 1874 Funcion 0.26375468
  when "011101010011"=> s <="101000011001"; -- Argumento 1875 Funcion 0.26227471
  when "011101010100"=> s <="101000010110"; -- Argumento 1876 Funcion 0.26079412
  when "011101010101"=> s <="101000010011"; -- Argumento 1877 Funcion 0.25931292
  when "011101010110"=> s <="101000010000"; -- Argumento 1878 Funcion 0.25783110
  when "011101010111"=> s <="101000001101"; -- Argumento 1879 Funcion 0.25634868
  when "011101011000"=> s <="101000001001"; -- Argumento 1880 Funcion 0.25486566
  when "011101011001"=> s <="101000000110"; -- Argumento 1881 Funcion 0.25338204
  when "011101011010"=> s <="101000000011"; -- Argumento 1882 Funcion 0.25189782
  when "011101011011"=> s <="101000000000"; -- Argumento 1883 Funcion 0.25041301
  when "011101011100"=> s <="100111111101"; -- Argumento 1884 Funcion 0.24892761
  when "011101011101"=> s <="100111111010"; -- Argumento 1885 Funcion 0.24744162
  when "011101011110"=> s <="100111110111"; -- Argumento 1886 Funcion 0.24595505
  when "011101011111"=> s <="100111110100"; -- Argumento 1887 Funcion 0.24446790
  when "011101100000"=> s <="100111110001"; -- Argumento 1888 Funcion 0.24298018
  when "011101100001"=> s <="100111101110"; -- Argumento 1889 Funcion 0.24149189
  when "011101100010"=> s <="100111101011"; -- Argumento 1890 Funcion 0.24000302
  when "011101100011"=> s <="100111101000"; -- Argumento 1891 Funcion 0.23851359
  when "011101100100"=> s <="100111100101"; -- Argumento 1892 Funcion 0.23702361
  when "011101100101"=> s <="100111100010"; -- Argumento 1893 Funcion 0.23553306
  when "011101100110"=> s <="100111011111"; -- Argumento 1894 Funcion 0.23404196
  when "011101100111"=> s <="100111011100"; -- Argumento 1895 Funcion 0.23255031
  when "011101101000"=> s <="100111011001"; -- Argumento 1896 Funcion 0.23105811
  when "011101101001"=> s <="100111010110"; -- Argumento 1897 Funcion 0.22956537
  when "011101101010"=> s <="100111010011"; -- Argumento 1898 Funcion 0.22807208
  when "011101101011"=> s <="100111010000"; -- Argumento 1899 Funcion 0.22657826
  when "011101101100"=> s <="100111001100"; -- Argumento 1900 Funcion 0.22508391
  when "011101101101"=> s <="100111001001"; -- Argumento 1901 Funcion 0.22358903
  when "011101101110"=> s <="100111000110"; -- Argumento 1902 Funcion 0.22209362
  when "011101101111"=> s <="100111000011"; -- Argumento 1903 Funcion 0.22059769
  when "011101110000"=> s <="100111000000"; -- Argumento 1904 Funcion 0.21910124
  when "011101110001"=> s <="100110111101"; -- Argumento 1905 Funcion 0.21760427
  when "011101110010"=> s <="100110111010"; -- Argumento 1906 Funcion 0.21610680
  when "011101110011"=> s <="100110110111"; -- Argumento 1907 Funcion 0.21460881
  when "011101110100"=> s <="100110110100"; -- Argumento 1908 Funcion 0.21311032
  when "011101110101"=> s <="100110110001"; -- Argumento 1909 Funcion 0.21161133
  when "011101110110"=> s <="100110101110"; -- Argumento 1910 Funcion 0.21011184
  when "011101110111"=> s <="100110101011"; -- Argumento 1911 Funcion 0.20861185
  when "011101111000"=> s <="100110101000"; -- Argumento 1912 Funcion 0.20711138
  when "011101111001"=> s <="100110100101"; -- Argumento 1913 Funcion 0.20561041
  when "011101111010"=> s <="100110100010"; -- Argumento 1914 Funcion 0.20410897
  when "011101111011"=> s <="100110011110"; -- Argumento 1915 Funcion 0.20260704
  when "011101111100"=> s <="100110011011"; -- Argumento 1916 Funcion 0.20110463
  when "011101111101"=> s <="100110011000"; -- Argumento 1917 Funcion 0.19960176
  when "011101111110"=> s <="100110010101"; -- Argumento 1918 Funcion 0.19809841
  when "011101111111"=> s <="100110010010"; -- Argumento 1919 Funcion 0.19659460
  when "011110000000"=> s <="100110001111"; -- Argumento 1920 Funcion 0.19509032
  when "011110000001"=> s <="100110001100"; -- Argumento 1921 Funcion 0.19358559
  when "011110000010"=> s <="100110001001"; -- Argumento 1922 Funcion 0.19208040
  when "011110000011"=> s <="100110000110"; -- Argumento 1923 Funcion 0.19057475
  when "011110000100"=> s <="100110000011"; -- Argumento 1924 Funcion 0.18906866
  when "011110000101"=> s <="100110000000"; -- Argumento 1925 Funcion 0.18756213
  when "011110000110"=> s <="100101111101"; -- Argumento 1926 Funcion 0.18605515
  when "011110000111"=> s <="100101111001"; -- Argumento 1927 Funcion 0.18454774
  when "011110001000"=> s <="100101110110"; -- Argumento 1928 Funcion 0.18303989
  when "011110001001"=> s <="100101110011"; -- Argumento 1929 Funcion 0.18153161
  when "011110001010"=> s <="100101110000"; -- Argumento 1930 Funcion 0.18002290
  when "011110001011"=> s <="100101101101"; -- Argumento 1931 Funcion 0.17851377
  when "011110001100"=> s <="100101101010"; -- Argumento 1932 Funcion 0.17700422
  when "011110001101"=> s <="100101100111"; -- Argumento 1933 Funcion 0.17549425
  when "011110001110"=> s <="100101100100"; -- Argumento 1934 Funcion 0.17398387
  when "011110001111"=> s <="100101100001"; -- Argumento 1935 Funcion 0.17247308
  when "011110010000"=> s <="100101011110"; -- Argumento 1936 Funcion 0.17096189
  when "011110010001"=> s <="100101011011"; -- Argumento 1937 Funcion 0.16945029
  when "011110010010"=> s <="100101010111"; -- Argumento 1938 Funcion 0.16793829
  when "011110010011"=> s <="100101010100"; -- Argumento 1939 Funcion 0.16642590
  when "011110010100"=> s <="100101010001"; -- Argumento 1940 Funcion 0.16491312
  when "011110010101"=> s <="100101001110"; -- Argumento 1941 Funcion 0.16339995
  when "011110010110"=> s <="100101001011"; -- Argumento 1942 Funcion 0.16188639
  when "011110010111"=> s <="100101001000"; -- Argumento 1943 Funcion 0.16037246
  when "011110011000"=> s <="100101000101"; -- Argumento 1944 Funcion 0.15885814
  when "011110011001"=> s <="100101000010"; -- Argumento 1945 Funcion 0.15734346
  when "011110011010"=> s <="100100111111"; -- Argumento 1946 Funcion 0.15582840
  when "011110011011"=> s <="100100111100"; -- Argumento 1947 Funcion 0.15431297
  when "011110011100"=> s <="100100111000"; -- Argumento 1948 Funcion 0.15279719
  when "011110011101"=> s <="100100110101"; -- Argumento 1949 Funcion 0.15128104
  when "011110011110"=> s <="100100110010"; -- Argumento 1950 Funcion 0.14976453
  when "011110011111"=> s <="100100101111"; -- Argumento 1951 Funcion 0.14824768
  when "011110100000"=> s <="100100101100"; -- Argumento 1952 Funcion 0.14673047
  when "011110100001"=> s <="100100101001"; -- Argumento 1953 Funcion 0.14521292
  when "011110100010"=> s <="100100100110"; -- Argumento 1954 Funcion 0.14369503
  when "011110100011"=> s <="100100100011"; -- Argumento 1955 Funcion 0.14217680
  when "011110100100"=> s <="100100100000"; -- Argumento 1956 Funcion 0.14065824
  when "011110100101"=> s <="100100011100"; -- Argumento 1957 Funcion 0.13913934
  when "011110100110"=> s <="100100011001"; -- Argumento 1958 Funcion 0.13762012
  when "011110100111"=> s <="100100010110"; -- Argumento 1959 Funcion 0.13610058
  when "011110101000"=> s <="100100010011"; -- Argumento 1960 Funcion 0.13458071
  when "011110101001"=> s <="100100010000"; -- Argumento 1961 Funcion 0.13306053
  when "011110101010"=> s <="100100001101"; -- Argumento 1962 Funcion 0.13154003
  when "011110101011"=> s <="100100001010"; -- Argumento 1963 Funcion 0.13001922
  when "011110101100"=> s <="100100000111"; -- Argumento 1964 Funcion 0.12849811
  when "011110101101"=> s <="100100000100"; -- Argumento 1965 Funcion 0.12697670
  when "011110101110"=> s <="100100000000"; -- Argumento 1966 Funcion 0.12545498
  when "011110101111"=> s <="100011111101"; -- Argumento 1967 Funcion 0.12393298
  when "011110110000"=> s <="100011111010"; -- Argumento 1968 Funcion 0.12241068
  when "011110110001"=> s <="100011110111"; -- Argumento 1969 Funcion 0.12088809
  when "011110110010"=> s <="100011110100"; -- Argumento 1970 Funcion 0.11936521
  when "011110110011"=> s <="100011110001"; -- Argumento 1971 Funcion 0.11784206
  when "011110110100"=> s <="100011101110"; -- Argumento 1972 Funcion 0.11631863
  when "011110110101"=> s <="100011101011"; -- Argumento 1973 Funcion 0.11479493
  when "011110110110"=> s <="100011100111"; -- Argumento 1974 Funcion 0.11327095
  when "011110110111"=> s <="100011100100"; -- Argumento 1975 Funcion 0.11174671
  when "011110111000"=> s <="100011100001"; -- Argumento 1976 Funcion 0.11022221
  when "011110111001"=> s <="100011011110"; -- Argumento 1977 Funcion 0.10869744
  when "011110111010"=> s <="100011011011"; -- Argumento 1978 Funcion 0.10717242
  when "011110111011"=> s <="100011011000"; -- Argumento 1979 Funcion 0.10564715
  when "011110111100"=> s <="100011010101"; -- Argumento 1980 Funcion 0.10412163
  when "011110111101"=> s <="100011010010"; -- Argumento 1981 Funcion 0.10259587
  when "011110111110"=> s <="100011001110"; -- Argumento 1982 Funcion 0.10106986
  when "011110111111"=> s <="100011001011"; -- Argumento 1983 Funcion 0.09954362
  when "011111000000"=> s <="100011001000"; -- Argumento 1984 Funcion 0.09801714
  when "011111000001"=> s <="100011000101"; -- Argumento 1985 Funcion 0.09649043
  when "011111000010"=> s <="100011000010"; -- Argumento 1986 Funcion 0.09496350
  when "011111000011"=> s <="100010111111"; -- Argumento 1987 Funcion 0.09343634
  when "011111000100"=> s <="100010111100"; -- Argumento 1988 Funcion 0.09190896
  when "011111000101"=> s <="100010111001"; -- Argumento 1989 Funcion 0.09038136
  when "011111000110"=> s <="100010110101"; -- Argumento 1990 Funcion 0.08885355
  when "011111000111"=> s <="100010110010"; -- Argumento 1991 Funcion 0.08732554
  when "011111001000"=> s <="100010101111"; -- Argumento 1992 Funcion 0.08579731
  when "011111001001"=> s <="100010101100"; -- Argumento 1993 Funcion 0.08426889
  when "011111001010"=> s <="100010101001"; -- Argumento 1994 Funcion 0.08274026
  when "011111001011"=> s <="100010100110"; -- Argumento 1995 Funcion 0.08121145
  when "011111001100"=> s <="100010100011"; -- Argumento 1996 Funcion 0.07968244
  when "011111001101"=> s <="100010100000"; -- Argumento 1997 Funcion 0.07815324
  when "011111001110"=> s <="100010011100"; -- Argumento 1998 Funcion 0.07662386
  when "011111001111"=> s <="100010011001"; -- Argumento 1999 Funcion 0.07509430
  when "011111010000"=> s <="100010010110"; -- Argumento 2000 Funcion 0.07356456
  when "011111010001"=> s <="100010010011"; -- Argumento 2001 Funcion 0.07203465
  when "011111010010"=> s <="100010010000"; -- Argumento 2002 Funcion 0.07050457
  when "011111010011"=> s <="100010001101"; -- Argumento 2003 Funcion 0.06897433
  when "011111010100"=> s <="100010001010"; -- Argumento 2004 Funcion 0.06744392
  when "011111010101"=> s <="100010000110"; -- Argumento 2005 Funcion 0.06591335
  when "011111010110"=> s <="100010000011"; -- Argumento 2006 Funcion 0.06438263
  when "011111010111"=> s <="100010000000"; -- Argumento 2007 Funcion 0.06285176
  when "011111011000"=> s <="100001111101"; -- Argumento 2008 Funcion 0.06132074
  when "011111011001"=> s <="100001111010"; -- Argumento 2009 Funcion 0.05978957
  when "011111011010"=> s <="100001110111"; -- Argumento 2010 Funcion 0.05825826
  when "011111011011"=> s <="100001110100"; -- Argumento 2011 Funcion 0.05672682
  when "011111011100"=> s <="100001110001"; -- Argumento 2012 Funcion 0.05519524
  when "011111011101"=> s <="100001101101"; -- Argumento 2013 Funcion 0.05366354
  when "011111011110"=> s <="100001101010"; -- Argumento 2014 Funcion 0.05213170
  when "011111011111"=> s <="100001100111"; -- Argumento 2015 Funcion 0.05059975
  when "011111100000"=> s <="100001100100"; -- Argumento 2016 Funcion 0.04906767
  when "011111100001"=> s <="100001100001"; -- Argumento 2017 Funcion 0.04753548
  when "011111100010"=> s <="100001011110"; -- Argumento 2018 Funcion 0.04600318
  when "011111100011"=> s <="100001011011"; -- Argumento 2019 Funcion 0.04447077
  when "011111100100"=> s <="100001010111"; -- Argumento 2020 Funcion 0.04293826
  when "011111100101"=> s <="100001010100"; -- Argumento 2021 Funcion 0.04140564
  when "011111100110"=> s <="100001010001"; -- Argumento 2022 Funcion 0.03987293
  when "011111100111"=> s <="100001001110"; -- Argumento 2023 Funcion 0.03834012
  when "011111101000"=> s <="100001001011"; -- Argumento 2024 Funcion 0.03680722
  when "011111101001"=> s <="100001001000"; -- Argumento 2025 Funcion 0.03527424
  when "011111101010"=> s <="100001000101"; -- Argumento 2026 Funcion 0.03374117
  when "011111101011"=> s <="100001000001"; -- Argumento 2027 Funcion 0.03220803
  when "011111101100"=> s <="100000111110"; -- Argumento 2028 Funcion 0.03067480
  when "011111101101"=> s <="100000111011"; -- Argumento 2029 Funcion 0.02914151
  when "011111101110"=> s <="100000111000"; -- Argumento 2030 Funcion 0.02760815
  when "011111101111"=> s <="100000110101"; -- Argumento 2031 Funcion 0.02607472
  when "011111110000"=> s <="100000110010"; -- Argumento 2032 Funcion 0.02454123
  when "011111110001"=> s <="100000101111"; -- Argumento 2033 Funcion 0.02300768
  when "011111110010"=> s <="100000101011"; -- Argumento 2034 Funcion 0.02147408
  when "011111110011"=> s <="100000101000"; -- Argumento 2035 Funcion 0.01994043
  when "011111110100"=> s <="100000100101"; -- Argumento 2036 Funcion 0.01840673
  when "011111110101"=> s <="100000100010"; -- Argumento 2037 Funcion 0.01687299
  when "011111110110"=> s <="100000011111"; -- Argumento 2038 Funcion 0.01533921
  when "011111110111"=> s <="100000011100"; -- Argumento 2039 Funcion 0.01380539
  when "011111111000"=> s <="100000011001"; -- Argumento 2040 Funcion 0.01227154
  when "011111111001"=> s <="100000010101"; -- Argumento 2041 Funcion 0.01073766
  when "011111111010"=> s <="100000010010"; -- Argumento 2042 Funcion 0.00920375
  when "011111111011"=> s <="100000001111"; -- Argumento 2043 Funcion 0.00766983
  when "011111111100"=> s <="100000001100"; -- Argumento 2044 Funcion 0.00613588
  when "011111111101"=> s <="100000001001"; -- Argumento 2045 Funcion 0.00460193
  when "011111111110"=> s <="100000000110"; -- Argumento 2046 Funcion 0.00306796
  when "011111111111"=> s <="100000000011"; -- Argumento 2047 Funcion 0.00153398
  when "100000000000"=> s <="100000000000"; -- Argumento 2048 Funcion 0.00000000
  when "100000000001"=> s <="011111111100"; -- Argumento 2049 Funcion -0.00153398
  when "100000000010"=> s <="011111111001"; -- Argumento 2050 Funcion -0.00306796
  when "100000000011"=> s <="011111110110"; -- Argumento 2051 Funcion -0.00460193
  when "100000000100"=> s <="011111110011"; -- Argumento 2052 Funcion -0.00613588
  when "100000000101"=> s <="011111110000"; -- Argumento 2053 Funcion -0.00766983
  when "100000000110"=> s <="011111101101"; -- Argumento 2054 Funcion -0.00920375
  when "100000000111"=> s <="011111101010"; -- Argumento 2055 Funcion -0.01073766
  when "100000001000"=> s <="011111100110"; -- Argumento 2056 Funcion -0.01227154
  when "100000001001"=> s <="011111100011"; -- Argumento 2057 Funcion -0.01380539
  when "100000001010"=> s <="011111100000"; -- Argumento 2058 Funcion -0.01533921
  when "100000001011"=> s <="011111011101"; -- Argumento 2059 Funcion -0.01687299
  when "100000001100"=> s <="011111011010"; -- Argumento 2060 Funcion -0.01840673
  when "100000001101"=> s <="011111010111"; -- Argumento 2061 Funcion -0.01994043
  when "100000001110"=> s <="011111010100"; -- Argumento 2062 Funcion -0.02147408
  when "100000001111"=> s <="011111010000"; -- Argumento 2063 Funcion -0.02300768
  when "100000010000"=> s <="011111001101"; -- Argumento 2064 Funcion -0.02454123
  when "100000010001"=> s <="011111001010"; -- Argumento 2065 Funcion -0.02607472
  when "100000010010"=> s <="011111000111"; -- Argumento 2066 Funcion -0.02760815
  when "100000010011"=> s <="011111000100"; -- Argumento 2067 Funcion -0.02914151
  when "100000010100"=> s <="011111000001"; -- Argumento 2068 Funcion -0.03067480
  when "100000010101"=> s <="011110111110"; -- Argumento 2069 Funcion -0.03220803
  when "100000010110"=> s <="011110111010"; -- Argumento 2070 Funcion -0.03374117
  when "100000010111"=> s <="011110110111"; -- Argumento 2071 Funcion -0.03527424
  when "100000011000"=> s <="011110110100"; -- Argumento 2072 Funcion -0.03680722
  when "100000011001"=> s <="011110110001"; -- Argumento 2073 Funcion -0.03834012
  when "100000011010"=> s <="011110101110"; -- Argumento 2074 Funcion -0.03987293
  when "100000011011"=> s <="011110101011"; -- Argumento 2075 Funcion -0.04140564
  when "100000011100"=> s <="011110101000"; -- Argumento 2076 Funcion -0.04293826
  when "100000011101"=> s <="011110100100"; -- Argumento 2077 Funcion -0.04447077
  when "100000011110"=> s <="011110100001"; -- Argumento 2078 Funcion -0.04600318
  when "100000011111"=> s <="011110011110"; -- Argumento 2079 Funcion -0.04753548
  when "100000100000"=> s <="011110011011"; -- Argumento 2080 Funcion -0.04906767
  when "100000100001"=> s <="011110011000"; -- Argumento 2081 Funcion -0.05059975
  when "100000100010"=> s <="011110010101"; -- Argumento 2082 Funcion -0.05213170
  when "100000100011"=> s <="011110010010"; -- Argumento 2083 Funcion -0.05366354
  when "100000100100"=> s <="011110001110"; -- Argumento 2084 Funcion -0.05519524
  when "100000100101"=> s <="011110001011"; -- Argumento 2085 Funcion -0.05672682
  when "100000100110"=> s <="011110001000"; -- Argumento 2086 Funcion -0.05825826
  when "100000100111"=> s <="011110000101"; -- Argumento 2087 Funcion -0.05978957
  when "100000101000"=> s <="011110000010"; -- Argumento 2088 Funcion -0.06132074
  when "100000101001"=> s <="011101111111"; -- Argumento 2089 Funcion -0.06285176
  when "100000101010"=> s <="011101111100"; -- Argumento 2090 Funcion -0.06438263
  when "100000101011"=> s <="011101111001"; -- Argumento 2091 Funcion -0.06591335
  when "100000101100"=> s <="011101110101"; -- Argumento 2092 Funcion -0.06744392
  when "100000101101"=> s <="011101110010"; -- Argumento 2093 Funcion -0.06897433
  when "100000101110"=> s <="011101101111"; -- Argumento 2094 Funcion -0.07050457
  when "100000101111"=> s <="011101101100"; -- Argumento 2095 Funcion -0.07203465
  when "100000110000"=> s <="011101101001"; -- Argumento 2096 Funcion -0.07356456
  when "100000110001"=> s <="011101100110"; -- Argumento 2097 Funcion -0.07509430
  when "100000110010"=> s <="011101100011"; -- Argumento 2098 Funcion -0.07662386
  when "100000110011"=> s <="011101011111"; -- Argumento 2099 Funcion -0.07815324
  when "100000110100"=> s <="011101011100"; -- Argumento 2100 Funcion -0.07968244
  when "100000110101"=> s <="011101011001"; -- Argumento 2101 Funcion -0.08121145
  when "100000110110"=> s <="011101010110"; -- Argumento 2102 Funcion -0.08274026
  when "100000110111"=> s <="011101010011"; -- Argumento 2103 Funcion -0.08426889
  when "100000111000"=> s <="011101010000"; -- Argumento 2104 Funcion -0.08579731
  when "100000111001"=> s <="011101001101"; -- Argumento 2105 Funcion -0.08732554
  when "100000111010"=> s <="011101001010"; -- Argumento 2106 Funcion -0.08885355
  when "100000111011"=> s <="011101000110"; -- Argumento 2107 Funcion -0.09038136
  when "100000111100"=> s <="011101000011"; -- Argumento 2108 Funcion -0.09190896
  when "100000111101"=> s <="011101000000"; -- Argumento 2109 Funcion -0.09343634
  when "100000111110"=> s <="011100111101"; -- Argumento 2110 Funcion -0.09496350
  when "100000111111"=> s <="011100111010"; -- Argumento 2111 Funcion -0.09649043
  when "100001000000"=> s <="011100110111"; -- Argumento 2112 Funcion -0.09801714
  when "100001000001"=> s <="011100110100"; -- Argumento 2113 Funcion -0.09954362
  when "100001000010"=> s <="011100110001"; -- Argumento 2114 Funcion -0.10106986
  when "100001000011"=> s <="011100101101"; -- Argumento 2115 Funcion -0.10259587
  when "100001000100"=> s <="011100101010"; -- Argumento 2116 Funcion -0.10412163
  when "100001000101"=> s <="011100100111"; -- Argumento 2117 Funcion -0.10564715
  when "100001000110"=> s <="011100100100"; -- Argumento 2118 Funcion -0.10717242
  when "100001000111"=> s <="011100100001"; -- Argumento 2119 Funcion -0.10869744
  when "100001001000"=> s <="011100011110"; -- Argumento 2120 Funcion -0.11022221
  when "100001001001"=> s <="011100011011"; -- Argumento 2121 Funcion -0.11174671
  when "100001001010"=> s <="011100011000"; -- Argumento 2122 Funcion -0.11327095
  when "100001001011"=> s <="011100010100"; -- Argumento 2123 Funcion -0.11479493
  when "100001001100"=> s <="011100010001"; -- Argumento 2124 Funcion -0.11631863
  when "100001001101"=> s <="011100001110"; -- Argumento 2125 Funcion -0.11784206
  when "100001001110"=> s <="011100001011"; -- Argumento 2126 Funcion -0.11936521
  when "100001001111"=> s <="011100001000"; -- Argumento 2127 Funcion -0.12088809
  when "100001010000"=> s <="011100000101"; -- Argumento 2128 Funcion -0.12241068
  when "100001010001"=> s <="011100000010"; -- Argumento 2129 Funcion -0.12393298
  when "100001010010"=> s <="011011111111"; -- Argumento 2130 Funcion -0.12545498
  when "100001010011"=> s <="011011111011"; -- Argumento 2131 Funcion -0.12697670
  when "100001010100"=> s <="011011111000"; -- Argumento 2132 Funcion -0.12849811
  when "100001010101"=> s <="011011110101"; -- Argumento 2133 Funcion -0.13001922
  when "100001010110"=> s <="011011110010"; -- Argumento 2134 Funcion -0.13154003
  when "100001010111"=> s <="011011101111"; -- Argumento 2135 Funcion -0.13306053
  when "100001011000"=> s <="011011101100"; -- Argumento 2136 Funcion -0.13458071
  when "100001011001"=> s <="011011101001"; -- Argumento 2137 Funcion -0.13610058
  when "100001011010"=> s <="011011100110"; -- Argumento 2138 Funcion -0.13762012
  when "100001011011"=> s <="011011100011"; -- Argumento 2139 Funcion -0.13913934
  when "100001011100"=> s <="011011011111"; -- Argumento 2140 Funcion -0.14065824
  when "100001011101"=> s <="011011011100"; -- Argumento 2141 Funcion -0.14217680
  when "100001011110"=> s <="011011011001"; -- Argumento 2142 Funcion -0.14369503
  when "100001011111"=> s <="011011010110"; -- Argumento 2143 Funcion -0.14521292
  when "100001100000"=> s <="011011010011"; -- Argumento 2144 Funcion -0.14673047
  when "100001100001"=> s <="011011010000"; -- Argumento 2145 Funcion -0.14824768
  when "100001100010"=> s <="011011001101"; -- Argumento 2146 Funcion -0.14976453
  when "100001100011"=> s <="011011001010"; -- Argumento 2147 Funcion -0.15128104
  when "100001100100"=> s <="011011000111"; -- Argumento 2148 Funcion -0.15279719
  when "100001100101"=> s <="011011000011"; -- Argumento 2149 Funcion -0.15431297
  when "100001100110"=> s <="011011000000"; -- Argumento 2150 Funcion -0.15582840
  when "100001100111"=> s <="011010111101"; -- Argumento 2151 Funcion -0.15734346
  when "100001101000"=> s <="011010111010"; -- Argumento 2152 Funcion -0.15885814
  when "100001101001"=> s <="011010110111"; -- Argumento 2153 Funcion -0.16037246
  when "100001101010"=> s <="011010110100"; -- Argumento 2154 Funcion -0.16188639
  when "100001101011"=> s <="011010110001"; -- Argumento 2155 Funcion -0.16339995
  when "100001101100"=> s <="011010101110"; -- Argumento 2156 Funcion -0.16491312
  when "100001101101"=> s <="011010101011"; -- Argumento 2157 Funcion -0.16642590
  when "100001101110"=> s <="011010101000"; -- Argumento 2158 Funcion -0.16793829
  when "100001101111"=> s <="011010100100"; -- Argumento 2159 Funcion -0.16945029
  when "100001110000"=> s <="011010100001"; -- Argumento 2160 Funcion -0.17096189
  when "100001110001"=> s <="011010011110"; -- Argumento 2161 Funcion -0.17247308
  when "100001110010"=> s <="011010011011"; -- Argumento 2162 Funcion -0.17398387
  when "100001110011"=> s <="011010011000"; -- Argumento 2163 Funcion -0.17549425
  when "100001110100"=> s <="011010010101"; -- Argumento 2164 Funcion -0.17700422
  when "100001110101"=> s <="011010010010"; -- Argumento 2165 Funcion -0.17851377
  when "100001110110"=> s <="011010001111"; -- Argumento 2166 Funcion -0.18002290
  when "100001110111"=> s <="011010001100"; -- Argumento 2167 Funcion -0.18153161
  when "100001111000"=> s <="011010001001"; -- Argumento 2168 Funcion -0.18303989
  when "100001111001"=> s <="011010000110"; -- Argumento 2169 Funcion -0.18454774
  when "100001111010"=> s <="011010000010"; -- Argumento 2170 Funcion -0.18605515
  when "100001111011"=> s <="011001111111"; -- Argumento 2171 Funcion -0.18756213
  when "100001111100"=> s <="011001111100"; -- Argumento 2172 Funcion -0.18906866
  when "100001111101"=> s <="011001111001"; -- Argumento 2173 Funcion -0.19057475
  when "100001111110"=> s <="011001110110"; -- Argumento 2174 Funcion -0.19208040
  when "100001111111"=> s <="011001110011"; -- Argumento 2175 Funcion -0.19358559
  when "100010000000"=> s <="011001110000"; -- Argumento 2176 Funcion -0.19509032
  when "100010000001"=> s <="011001101101"; -- Argumento 2177 Funcion -0.19659460
  when "100010000010"=> s <="011001101010"; -- Argumento 2178 Funcion -0.19809841
  when "100010000011"=> s <="011001100111"; -- Argumento 2179 Funcion -0.19960176
  when "100010000100"=> s <="011001100100"; -- Argumento 2180 Funcion -0.20110463
  when "100010000101"=> s <="011001100001"; -- Argumento 2181 Funcion -0.20260704
  when "100010000110"=> s <="011001011101"; -- Argumento 2182 Funcion -0.20410897
  when "100010000111"=> s <="011001011010"; -- Argumento 2183 Funcion -0.20561041
  when "100010001000"=> s <="011001010111"; -- Argumento 2184 Funcion -0.20711138
  when "100010001001"=> s <="011001010100"; -- Argumento 2185 Funcion -0.20861185
  when "100010001010"=> s <="011001010001"; -- Argumento 2186 Funcion -0.21011184
  when "100010001011"=> s <="011001001110"; -- Argumento 2187 Funcion -0.21161133
  when "100010001100"=> s <="011001001011"; -- Argumento 2188 Funcion -0.21311032
  when "100010001101"=> s <="011001001000"; -- Argumento 2189 Funcion -0.21460881
  when "100010001110"=> s <="011001000101"; -- Argumento 2190 Funcion -0.21610680
  when "100010001111"=> s <="011001000010"; -- Argumento 2191 Funcion -0.21760427
  when "100010010000"=> s <="011000111111"; -- Argumento 2192 Funcion -0.21910124
  when "100010010001"=> s <="011000111100"; -- Argumento 2193 Funcion -0.22059769
  when "100010010010"=> s <="011000111001"; -- Argumento 2194 Funcion -0.22209362
  when "100010010011"=> s <="011000110110"; -- Argumento 2195 Funcion -0.22358903
  when "100010010100"=> s <="011000110011"; -- Argumento 2196 Funcion -0.22508391
  when "100010010101"=> s <="011000101111"; -- Argumento 2197 Funcion -0.22657826
  when "100010010110"=> s <="011000101100"; -- Argumento 2198 Funcion -0.22807208
  when "100010010111"=> s <="011000101001"; -- Argumento 2199 Funcion -0.22956537
  when "100010011000"=> s <="011000100110"; -- Argumento 2200 Funcion -0.23105811
  when "100010011001"=> s <="011000100011"; -- Argumento 2201 Funcion -0.23255031
  when "100010011010"=> s <="011000100000"; -- Argumento 2202 Funcion -0.23404196
  when "100010011011"=> s <="011000011101"; -- Argumento 2203 Funcion -0.23553306
  when "100010011100"=> s <="011000011010"; -- Argumento 2204 Funcion -0.23702361
  when "100010011101"=> s <="011000010111"; -- Argumento 2205 Funcion -0.23851359
  when "100010011110"=> s <="011000010100"; -- Argumento 2206 Funcion -0.24000302
  when "100010011111"=> s <="011000010001"; -- Argumento 2207 Funcion -0.24149189
  when "100010100000"=> s <="011000001110"; -- Argumento 2208 Funcion -0.24298018
  when "100010100001"=> s <="011000001011"; -- Argumento 2209 Funcion -0.24446790
  when "100010100010"=> s <="011000001000"; -- Argumento 2210 Funcion -0.24595505
  when "100010100011"=> s <="011000000101"; -- Argumento 2211 Funcion -0.24744162
  when "100010100100"=> s <="011000000010"; -- Argumento 2212 Funcion -0.24892761
  when "100010100101"=> s <="010111111111"; -- Argumento 2213 Funcion -0.25041301
  when "100010100110"=> s <="010111111100"; -- Argumento 2214 Funcion -0.25189782
  when "100010100111"=> s <="010111111001"; -- Argumento 2215 Funcion -0.25338204
  when "100010101000"=> s <="010111110110"; -- Argumento 2216 Funcion -0.25486566
  when "100010101001"=> s <="010111110010"; -- Argumento 2217 Funcion -0.25634868
  when "100010101010"=> s <="010111101111"; -- Argumento 2218 Funcion -0.25783110
  when "100010101011"=> s <="010111101100"; -- Argumento 2219 Funcion -0.25931292
  when "100010101100"=> s <="010111101001"; -- Argumento 2220 Funcion -0.26079412
  when "100010101101"=> s <="010111100110"; -- Argumento 2221 Funcion -0.26227471
  when "100010101110"=> s <="010111100011"; -- Argumento 2222 Funcion -0.26375468
  when "100010101111"=> s <="010111100000"; -- Argumento 2223 Funcion -0.26523403
  when "100010110000"=> s <="010111011101"; -- Argumento 2224 Funcion -0.26671276
  when "100010110001"=> s <="010111011010"; -- Argumento 2225 Funcion -0.26819086
  when "100010110010"=> s <="010111010111"; -- Argumento 2226 Funcion -0.26966833
  when "100010110011"=> s <="010111010100"; -- Argumento 2227 Funcion -0.27114516
  when "100010110100"=> s <="010111010001"; -- Argumento 2228 Funcion -0.27262136
  when "100010110101"=> s <="010111001110"; -- Argumento 2229 Funcion -0.27409691
  when "100010110110"=> s <="010111001011"; -- Argumento 2230 Funcion -0.27557182
  when "100010110111"=> s <="010111001000"; -- Argumento 2231 Funcion -0.27704608
  when "100010111000"=> s <="010111000101"; -- Argumento 2232 Funcion -0.27851969
  when "100010111001"=> s <="010111000010"; -- Argumento 2233 Funcion -0.27999264
  when "100010111010"=> s <="010110111111"; -- Argumento 2234 Funcion -0.28146494
  when "100010111011"=> s <="010110111100"; -- Argumento 2235 Funcion -0.28293657
  when "100010111100"=> s <="010110111001"; -- Argumento 2236 Funcion -0.28440754
  when "100010111101"=> s <="010110110110"; -- Argumento 2237 Funcion -0.28587783
  when "100010111110"=> s <="010110110011"; -- Argumento 2238 Funcion -0.28734746
  when "100010111111"=> s <="010110110000"; -- Argumento 2239 Funcion -0.28881641
  when "100011000000"=> s <="010110101101"; -- Argumento 2240 Funcion -0.29028468
  when "100011000001"=> s <="010110101010"; -- Argumento 2241 Funcion -0.29175226
  when "100011000010"=> s <="010110100111"; -- Argumento 2242 Funcion -0.29321916
  when "100011000011"=> s <="010110100100"; -- Argumento 2243 Funcion -0.29468537
  when "100011000100"=> s <="010110100001"; -- Argumento 2244 Funcion -0.29615089
  when "100011000101"=> s <="010110011110"; -- Argumento 2245 Funcion -0.29761571
  when "100011000110"=> s <="010110011011"; -- Argumento 2246 Funcion -0.29907983
  when "100011000111"=> s <="010110011000"; -- Argumento 2247 Funcion -0.30054324
  when "100011001000"=> s <="010110010101"; -- Argumento 2248 Funcion -0.30200595
  when "100011001001"=> s <="010110010010"; -- Argumento 2249 Funcion -0.30346795
  when "100011001010"=> s <="010110001111"; -- Argumento 2250 Funcion -0.30492923
  when "100011001011"=> s <="010110001100"; -- Argumento 2251 Funcion -0.30638980
  when "100011001100"=> s <="010110001001"; -- Argumento 2252 Funcion -0.30784964
  when "100011001101"=> s <="010110000110"; -- Argumento 2253 Funcion -0.30930876
  when "100011001110"=> s <="010110000011"; -- Argumento 2254 Funcion -0.31076715
  when "100011001111"=> s <="010110000000"; -- Argumento 2255 Funcion -0.31222481
  when "100011010000"=> s <="010101111101"; -- Argumento 2256 Funcion -0.31368174
  when "100011010001"=> s <="010101111010"; -- Argumento 2257 Funcion -0.31513793
  when "100011010010"=> s <="010101110111"; -- Argumento 2258 Funcion -0.31659338
  when "100011010011"=> s <="010101110100"; -- Argumento 2259 Funcion -0.31804808
  when "100011010100"=> s <="010101110001"; -- Argumento 2260 Funcion -0.31950203
  when "100011010101"=> s <="010101101110"; -- Argumento 2261 Funcion -0.32095523
  when "100011010110"=> s <="010101101011"; -- Argumento 2262 Funcion -0.32240768
  when "100011010111"=> s <="010101101000"; -- Argumento 2263 Funcion -0.32385937
  when "100011011000"=> s <="010101100101"; -- Argumento 2264 Funcion -0.32531029
  when "100011011001"=> s <="010101100010"; -- Argumento 2265 Funcion -0.32676045
  when "100011011010"=> s <="010101011111"; -- Argumento 2266 Funcion -0.32820984
  when "100011011011"=> s <="010101011100"; -- Argumento 2267 Funcion -0.32965846
  when "100011011100"=> s <="010101011001"; -- Argumento 2268 Funcion -0.33110631
  when "100011011101"=> s <="010101010110"; -- Argumento 2269 Funcion -0.33255337
  when "100011011110"=> s <="010101010011"; -- Argumento 2270 Funcion -0.33399965
  when "100011011111"=> s <="010101010001"; -- Argumento 2271 Funcion -0.33544515
  when "100011100000"=> s <="010101001110"; -- Argumento 2272 Funcion -0.33688985
  when "100011100001"=> s <="010101001011"; -- Argumento 2273 Funcion -0.33833377
  when "100011100010"=> s <="010101001000"; -- Argumento 2274 Funcion -0.33977688
  when "100011100011"=> s <="010101000101"; -- Argumento 2275 Funcion -0.34121920
  when "100011100100"=> s <="010101000010"; -- Argumento 2276 Funcion -0.34266072
  when "100011100101"=> s <="010100111111"; -- Argumento 2277 Funcion -0.34410143
  when "100011100110"=> s <="010100111100"; -- Argumento 2278 Funcion -0.34554132
  when "100011100111"=> s <="010100111001"; -- Argumento 2279 Funcion -0.34698041
  when "100011101000"=> s <="010100110110"; -- Argumento 2280 Funcion -0.34841868
  when "100011101001"=> s <="010100110011"; -- Argumento 2281 Funcion -0.34985613
  when "100011101010"=> s <="010100110000"; -- Argumento 2282 Funcion -0.35129276
  when "100011101011"=> s <="010100101101"; -- Argumento 2283 Funcion -0.35272856
  when "100011101100"=> s <="010100101010"; -- Argumento 2284 Funcion -0.35416353
  when "100011101101"=> s <="010100100111"; -- Argumento 2285 Funcion -0.35559766
  when "100011101110"=> s <="010100100100"; -- Argumento 2286 Funcion -0.35703096
  when "100011101111"=> s <="010100100001"; -- Argumento 2287 Funcion -0.35846342
  when "100011110000"=> s <="010100011110"; -- Argumento 2288 Funcion -0.35989504
  when "100011110001"=> s <="010100011100"; -- Argumento 2289 Funcion -0.36132581
  when "100011110010"=> s <="010100011001"; -- Argumento 2290 Funcion -0.36275572
  when "100011110011"=> s <="010100010110"; -- Argumento 2291 Funcion -0.36418479
  when "100011110100"=> s <="010100010011"; -- Argumento 2292 Funcion -0.36561300
  when "100011110101"=> s <="010100010000"; -- Argumento 2293 Funcion -0.36704035
  when "100011110110"=> s <="010100001101"; -- Argumento 2294 Funcion -0.36846683
  when "100011110111"=> s <="010100001010"; -- Argumento 2295 Funcion -0.36989245
  when "100011111000"=> s <="010100000111"; -- Argumento 2296 Funcion -0.37131719
  when "100011111001"=> s <="010100000100"; -- Argumento 2297 Funcion -0.37274107
  when "100011111010"=> s <="010100000001"; -- Argumento 2298 Funcion -0.37416406
  when "100011111011"=> s <="010011111110"; -- Argumento 2299 Funcion -0.37558618
  when "100011111100"=> s <="010011111011"; -- Argumento 2300 Funcion -0.37700741
  when "100011111101"=> s <="010011111000"; -- Argumento 2301 Funcion -0.37842775
  when "100011111110"=> s <="010011110110"; -- Argumento 2302 Funcion -0.37984721
  when "100011111111"=> s <="010011110011"; -- Argumento 2303 Funcion -0.38126577
  when "100100000000"=> s <="010011110000"; -- Argumento 2304 Funcion -0.38268343
  when "100100000001"=> s <="010011101101"; -- Argumento 2305 Funcion -0.38410020
  when "100100000010"=> s <="010011101010"; -- Argumento 2306 Funcion -0.38551605
  when "100100000011"=> s <="010011100111"; -- Argumento 2307 Funcion -0.38693101
  when "100100000100"=> s <="010011100100"; -- Argumento 2308 Funcion -0.38834505
  when "100100000101"=> s <="010011100001"; -- Argumento 2309 Funcion -0.38975817
  when "100100000110"=> s <="010011011110"; -- Argumento 2310 Funcion -0.39117038
  when "100100000111"=> s <="010011011011"; -- Argumento 2311 Funcion -0.39258167
  when "100100001000"=> s <="010011011001"; -- Argumento 2312 Funcion -0.39399204
  when "100100001001"=> s <="010011010110"; -- Argumento 2313 Funcion -0.39540148
  when "100100001010"=> s <="010011010011"; -- Argumento 2314 Funcion -0.39680999
  when "100100001011"=> s <="010011010000"; -- Argumento 2315 Funcion -0.39821756
  when "100100001100"=> s <="010011001101"; -- Argumento 2316 Funcion -0.39962420
  when "100100001101"=> s <="010011001010"; -- Argumento 2317 Funcion -0.40102990
  when "100100001110"=> s <="010011000111"; -- Argumento 2318 Funcion -0.40243465
  when "100100001111"=> s <="010011000100"; -- Argumento 2319 Funcion -0.40383846
  when "100100010000"=> s <="010011000010"; -- Argumento 2320 Funcion -0.40524131
  when "100100010001"=> s <="010010111111"; -- Argumento 2321 Funcion -0.40664322
  when "100100010010"=> s <="010010111100"; -- Argumento 2322 Funcion -0.40804416
  when "100100010011"=> s <="010010111001"; -- Argumento 2323 Funcion -0.40944415
  when "100100010100"=> s <="010010110110"; -- Argumento 2324 Funcion -0.41084317
  when "100100010101"=> s <="010010110011"; -- Argumento 2325 Funcion -0.41224123
  when "100100010110"=> s <="010010110000"; -- Argumento 2326 Funcion -0.41363831
  when "100100010111"=> s <="010010101110"; -- Argumento 2327 Funcion -0.41503442
  when "100100011000"=> s <="010010101011"; -- Argumento 2328 Funcion -0.41642956
  when "100100011001"=> s <="010010101000"; -- Argumento 2329 Funcion -0.41782372
  when "100100011010"=> s <="010010100101"; -- Argumento 2330 Funcion -0.41921689
  when "100100011011"=> s <="010010100010"; -- Argumento 2331 Funcion -0.42060907
  when "100100011100"=> s <="010010011111"; -- Argumento 2332 Funcion -0.42200027
  when "100100011101"=> s <="010010011100"; -- Argumento 2333 Funcion -0.42339047
  when "100100011110"=> s <="010010011010"; -- Argumento 2334 Funcion -0.42477968
  when "100100011111"=> s <="010010010111"; -- Argumento 2335 Funcion -0.42616789
  when "100100100000"=> s <="010010010100"; -- Argumento 2336 Funcion -0.42755509
  when "100100100001"=> s <="010010010001"; -- Argumento 2337 Funcion -0.42894129
  when "100100100010"=> s <="010010001110"; -- Argumento 2338 Funcion -0.43032648
  when "100100100011"=> s <="010010001011"; -- Argumento 2339 Funcion -0.43171066
  when "100100100100"=> s <="010010001001"; -- Argumento 2340 Funcion -0.43309382
  when "100100100101"=> s <="010010000110"; -- Argumento 2341 Funcion -0.43447596
  when "100100100110"=> s <="010010000011"; -- Argumento 2342 Funcion -0.43585708
  when "100100100111"=> s <="010010000000"; -- Argumento 2343 Funcion -0.43723717
  when "100100101000"=> s <="010001111101"; -- Argumento 2344 Funcion -0.43861624
  when "100100101001"=> s <="010001111010"; -- Argumento 2345 Funcion -0.43999427
  when "100100101010"=> s <="010001111000"; -- Argumento 2346 Funcion -0.44137127
  when "100100101011"=> s <="010001110101"; -- Argumento 2347 Funcion -0.44274723
  when "100100101100"=> s <="010001110010"; -- Argumento 2348 Funcion -0.44412214
  when "100100101101"=> s <="010001101111"; -- Argumento 2349 Funcion -0.44549602
  when "100100101110"=> s <="010001101100"; -- Argumento 2350 Funcion -0.44686884
  when "100100101111"=> s <="010001101010"; -- Argumento 2351 Funcion -0.44824061
  when "100100110000"=> s <="010001100111"; -- Argumento 2352 Funcion -0.44961133
  when "100100110001"=> s <="010001100100"; -- Argumento 2353 Funcion -0.45098099
  when "100100110010"=> s <="010001100001"; -- Argumento 2354 Funcion -0.45234959
  when "100100110011"=> s <="010001011110"; -- Argumento 2355 Funcion -0.45371712
  when "100100110100"=> s <="010001011011"; -- Argumento 2356 Funcion -0.45508359
  when "100100110101"=> s <="010001011001"; -- Argumento 2357 Funcion -0.45644898
  when "100100110110"=> s <="010001010110"; -- Argumento 2358 Funcion -0.45781330
  when "100100110111"=> s <="010001010011"; -- Argumento 2359 Funcion -0.45917655
  when "100100111000"=> s <="010001010000"; -- Argumento 2360 Funcion -0.46053871
  when "100100111001"=> s <="010001001110"; -- Argumento 2361 Funcion -0.46189979
  when "100100111010"=> s <="010001001011"; -- Argumento 2362 Funcion -0.46325978
  when "100100111011"=> s <="010001001000"; -- Argumento 2363 Funcion -0.46461869
  when "100100111100"=> s <="010001000101"; -- Argumento 2364 Funcion -0.46597650
  when "100100111101"=> s <="010001000010"; -- Argumento 2365 Funcion -0.46733321
  when "100100111110"=> s <="010001000000"; -- Argumento 2366 Funcion -0.46868882
  when "100100111111"=> s <="010000111101"; -- Argumento 2367 Funcion -0.47004333
  when "100101000000"=> s <="010000111010"; -- Argumento 2368 Funcion -0.47139674
  when "100101000001"=> s <="010000110111"; -- Argumento 2369 Funcion -0.47274903
  when "100101000010"=> s <="010000110101"; -- Argumento 2370 Funcion -0.47410021
  when "100101000011"=> s <="010000110010"; -- Argumento 2371 Funcion -0.47545028
  when "100101000100"=> s <="010000101111"; -- Argumento 2372 Funcion -0.47679923
  when "100101000101"=> s <="010000101100"; -- Argumento 2373 Funcion -0.47814706
  when "100101000110"=> s <="010000101001"; -- Argumento 2374 Funcion -0.47949376
  when "100101000111"=> s <="010000100111"; -- Argumento 2375 Funcion -0.48083933
  when "100101001000"=> s <="010000100100"; -- Argumento 2376 Funcion -0.48218377
  when "100101001001"=> s <="010000100001"; -- Argumento 2377 Funcion -0.48352708
  when "100101001010"=> s <="010000011110"; -- Argumento 2378 Funcion -0.48486925
  when "100101001011"=> s <="010000011100"; -- Argumento 2379 Funcion -0.48621028
  when "100101001100"=> s <="010000011001"; -- Argumento 2380 Funcion -0.48755016
  when "100101001101"=> s <="010000010110"; -- Argumento 2381 Funcion -0.48888890
  when "100101001110"=> s <="010000010100"; -- Argumento 2382 Funcion -0.49022648
  when "100101001111"=> s <="010000010001"; -- Argumento 2383 Funcion -0.49156292
  when "100101010000"=> s <="010000001110"; -- Argumento 2384 Funcion -0.49289819
  when "100101010001"=> s <="010000001011"; -- Argumento 2385 Funcion -0.49423231
  when "100101010010"=> s <="010000001001"; -- Argumento 2386 Funcion -0.49556526
  when "100101010011"=> s <="010000000110"; -- Argumento 2387 Funcion -0.49689705
  when "100101010100"=> s <="010000000011"; -- Argumento 2388 Funcion -0.49822767
  when "100101010101"=> s <="010000000000"; -- Argumento 2389 Funcion -0.49955711
  when "100101010110"=> s <="001111111110"; -- Argumento 2390 Funcion -0.50088538
  when "100101010111"=> s <="001111111011"; -- Argumento 2391 Funcion -0.50221247
  when "100101011000"=> s <="001111111000"; -- Argumento 2392 Funcion -0.50353838
  when "100101011001"=> s <="001111110110"; -- Argumento 2393 Funcion -0.50486311
  when "100101011010"=> s <="001111110011"; -- Argumento 2394 Funcion -0.50618665
  when "100101011011"=> s <="001111110000"; -- Argumento 2395 Funcion -0.50750899
  when "100101011100"=> s <="001111101101"; -- Argumento 2396 Funcion -0.50883014
  when "100101011101"=> s <="001111101011"; -- Argumento 2397 Funcion -0.51015010
  when "100101011110"=> s <="001111101000"; -- Argumento 2398 Funcion -0.51146885
  when "100101011111"=> s <="001111100101"; -- Argumento 2399 Funcion -0.51278640
  when "100101100000"=> s <="001111100011"; -- Argumento 2400 Funcion -0.51410274
  when "100101100001"=> s <="001111100000"; -- Argumento 2401 Funcion -0.51541788
  when "100101100010"=> s <="001111011101"; -- Argumento 2402 Funcion -0.51673180
  when "100101100011"=> s <="001111011011"; -- Argumento 2403 Funcion -0.51804450
  when "100101100100"=> s <="001111011000"; -- Argumento 2404 Funcion -0.51935599
  when "100101100101"=> s <="001111010101"; -- Argumento 2405 Funcion -0.52066625
  when "100101100110"=> s <="001111010010"; -- Argumento 2406 Funcion -0.52197529
  when "100101100111"=> s <="001111010000"; -- Argumento 2407 Funcion -0.52328310
  when "100101101000"=> s <="001111001101"; -- Argumento 2408 Funcion -0.52458968
  when "100101101001"=> s <="001111001010"; -- Argumento 2409 Funcion -0.52589503
  when "100101101010"=> s <="001111001000"; -- Argumento 2410 Funcion -0.52719913
  when "100101101011"=> s <="001111000101"; -- Argumento 2411 Funcion -0.52850200
  when "100101101100"=> s <="001111000010"; -- Argumento 2412 Funcion -0.52980362
  when "100101101101"=> s <="001111000000"; -- Argumento 2413 Funcion -0.53110400
  when "100101101110"=> s <="001110111101"; -- Argumento 2414 Funcion -0.53240313
  when "100101101111"=> s <="001110111010"; -- Argumento 2415 Funcion -0.53370100
  when "100101110000"=> s <="001110111000"; -- Argumento 2416 Funcion -0.53499762
  when "100101110001"=> s <="001110110101"; -- Argumento 2417 Funcion -0.53629298
  when "100101110010"=> s <="001110110011"; -- Argumento 2418 Funcion -0.53758708
  when "100101110011"=> s <="001110110000"; -- Argumento 2419 Funcion -0.53887991
  when "100101110100"=> s <="001110101101"; -- Argumento 2420 Funcion -0.54017147
  when "100101110101"=> s <="001110101011"; -- Argumento 2421 Funcion -0.54146177
  when "100101110110"=> s <="001110101000"; -- Argumento 2422 Funcion -0.54275078
  when "100101110111"=> s <="001110100101"; -- Argumento 2423 Funcion -0.54403853
  when "100101111000"=> s <="001110100011"; -- Argumento 2424 Funcion -0.54532499
  when "100101111001"=> s <="001110100000"; -- Argumento 2425 Funcion -0.54661017
  when "100101111010"=> s <="001110011101"; -- Argumento 2426 Funcion -0.54789406
  when "100101111011"=> s <="001110011011"; -- Argumento 2427 Funcion -0.54917666
  when "100101111100"=> s <="001110011000"; -- Argumento 2428 Funcion -0.55045797
  when "100101111101"=> s <="001110010110"; -- Argumento 2429 Funcion -0.55173799
  when "100101111110"=> s <="001110010011"; -- Argumento 2430 Funcion -0.55301671
  when "100101111111"=> s <="001110010000"; -- Argumento 2431 Funcion -0.55429412
  when "100110000000"=> s <="001110001110"; -- Argumento 2432 Funcion -0.55557023
  when "100110000001"=> s <="001110001011"; -- Argumento 2433 Funcion -0.55684504
  when "100110000010"=> s <="001110001000"; -- Argumento 2434 Funcion -0.55811853
  when "100110000011"=> s <="001110000110"; -- Argumento 2435 Funcion -0.55939071
  when "100110000100"=> s <="001110000011"; -- Argumento 2436 Funcion -0.56066158
  when "100110000101"=> s <="001110000001"; -- Argumento 2437 Funcion -0.56193112
  when "100110000110"=> s <="001101111110"; -- Argumento 2438 Funcion -0.56319934
  when "100110000111"=> s <="001101111011"; -- Argumento 2439 Funcion -0.56446624
  when "100110001000"=> s <="001101111001"; -- Argumento 2440 Funcion -0.56573181
  when "100110001001"=> s <="001101110110"; -- Argumento 2441 Funcion -0.56699605
  when "100110001010"=> s <="001101110100"; -- Argumento 2442 Funcion -0.56825895
  when "100110001011"=> s <="001101110001"; -- Argumento 2443 Funcion -0.56952052
  when "100110001100"=> s <="001101101111"; -- Argumento 2444 Funcion -0.57078075
  when "100110001101"=> s <="001101101100"; -- Argumento 2445 Funcion -0.57203963
  when "100110001110"=> s <="001101101001"; -- Argumento 2446 Funcion -0.57329717
  when "100110001111"=> s <="001101100111"; -- Argumento 2447 Funcion -0.57455336
  when "100110010000"=> s <="001101100100"; -- Argumento 2448 Funcion -0.57580819
  when "100110010001"=> s <="001101100010"; -- Argumento 2449 Funcion -0.57706167
  when "100110010010"=> s <="001101011111"; -- Argumento 2450 Funcion -0.57831380
  when "100110010011"=> s <="001101011101"; -- Argumento 2451 Funcion -0.57956456
  when "100110010100"=> s <="001101011010"; -- Argumento 2452 Funcion -0.58081396
  when "100110010101"=> s <="001101010111"; -- Argumento 2453 Funcion -0.58206199
  when "100110010110"=> s <="001101010101"; -- Argumento 2454 Funcion -0.58330865
  when "100110010111"=> s <="001101010010"; -- Argumento 2455 Funcion -0.58455394
  when "100110011000"=> s <="001101010000"; -- Argumento 2456 Funcion -0.58579786
  when "100110011001"=> s <="001101001101"; -- Argumento 2457 Funcion -0.58704039
  when "100110011010"=> s <="001101001011"; -- Argumento 2458 Funcion -0.58828155
  when "100110011011"=> s <="001101001000"; -- Argumento 2459 Funcion -0.58952132
  when "100110011100"=> s <="001101000110"; -- Argumento 2460 Funcion -0.59075970
  when "100110011101"=> s <="001101000011"; -- Argumento 2461 Funcion -0.59199669
  when "100110011110"=> s <="001101000001"; -- Argumento 2462 Funcion -0.59323230
  when "100110011111"=> s <="001100111110"; -- Argumento 2463 Funcion -0.59446650
  when "100110100000"=> s <="001100111100"; -- Argumento 2464 Funcion -0.59569930
  when "100110100001"=> s <="001100111001"; -- Argumento 2465 Funcion -0.59693071
  when "100110100010"=> s <="001100110110"; -- Argumento 2466 Funcion -0.59816071
  when "100110100011"=> s <="001100110100"; -- Argumento 2467 Funcion -0.59938930
  when "100110100100"=> s <="001100110001"; -- Argumento 2468 Funcion -0.60061648
  when "100110100101"=> s <="001100101111"; -- Argumento 2469 Funcion -0.60184225
  when "100110100110"=> s <="001100101100"; -- Argumento 2470 Funcion -0.60306660
  when "100110100111"=> s <="001100101010"; -- Argumento 2471 Funcion -0.60428953
  when "100110101000"=> s <="001100100111"; -- Argumento 2472 Funcion -0.60551104
  when "100110101001"=> s <="001100100101"; -- Argumento 2473 Funcion -0.60673113
  when "100110101010"=> s <="001100100010"; -- Argumento 2474 Funcion -0.60794978
  when "100110101011"=> s <="001100100000"; -- Argumento 2475 Funcion -0.60916701
  when "100110101100"=> s <="001100011101"; -- Argumento 2476 Funcion -0.61038281
  when "100110101101"=> s <="001100011011"; -- Argumento 2477 Funcion -0.61159716
  when "100110101110"=> s <="001100011000"; -- Argumento 2478 Funcion -0.61281008
  when "100110101111"=> s <="001100010110"; -- Argumento 2479 Funcion -0.61402156
  when "100110110000"=> s <="001100010100"; -- Argumento 2480 Funcion -0.61523159
  when "100110110001"=> s <="001100010001"; -- Argumento 2481 Funcion -0.61644017
  when "100110110010"=> s <="001100001111"; -- Argumento 2482 Funcion -0.61764731
  when "100110110011"=> s <="001100001100"; -- Argumento 2483 Funcion -0.61885299
  when "100110110100"=> s <="001100001010"; -- Argumento 2484 Funcion -0.62005721
  when "100110110101"=> s <="001100000111"; -- Argumento 2485 Funcion -0.62125998
  when "100110110110"=> s <="001100000101"; -- Argumento 2486 Funcion -0.62246128
  when "100110110111"=> s <="001100000010"; -- Argumento 2487 Funcion -0.62366112
  when "100110111000"=> s <="001100000000"; -- Argumento 2488 Funcion -0.62485949
  when "100110111001"=> s <="001011111101"; -- Argumento 2489 Funcion -0.62605639
  when "100110111010"=> s <="001011111011"; -- Argumento 2490 Funcion -0.62725182
  when "100110111011"=> s <="001011111000"; -- Argumento 2491 Funcion -0.62844577
  when "100110111100"=> s <="001011110110"; -- Argumento 2492 Funcion -0.62963824
  when "100110111101"=> s <="001011110100"; -- Argumento 2493 Funcion -0.63082923
  when "100110111110"=> s <="001011110001"; -- Argumento 2494 Funcion -0.63201874
  when "100110111111"=> s <="001011101111"; -- Argumento 2495 Funcion -0.63320676
  when "100111000000"=> s <="001011101100"; -- Argumento 2496 Funcion -0.63439328
  when "100111000001"=> s <="001011101010"; -- Argumento 2497 Funcion -0.63557832
  when "100111000010"=> s <="001011100111"; -- Argumento 2498 Funcion -0.63676186
  when "100111000011"=> s <="001011100101"; -- Argumento 2499 Funcion -0.63794390
  when "100111000100"=> s <="001011100011"; -- Argumento 2500 Funcion -0.63912444
  when "100111000101"=> s <="001011100000"; -- Argumento 2501 Funcion -0.64030348
  when "100111000110"=> s <="001011011110"; -- Argumento 2502 Funcion -0.64148101
  when "100111000111"=> s <="001011011011"; -- Argumento 2503 Funcion -0.64265703
  when "100111001000"=> s <="001011011001"; -- Argumento 2504 Funcion -0.64383154
  when "100111001001"=> s <="001011010111"; -- Argumento 2505 Funcion -0.64500454
  when "100111001010"=> s <="001011010100"; -- Argumento 2506 Funcion -0.64617601
  when "100111001011"=> s <="001011010010"; -- Argumento 2507 Funcion -0.64734597
  when "100111001100"=> s <="001011001111"; -- Argumento 2508 Funcion -0.64851440
  when "100111001101"=> s <="001011001101"; -- Argumento 2509 Funcion -0.64968131
  when "100111001110"=> s <="001011001011"; -- Argumento 2510 Funcion -0.65084668
  when "100111001111"=> s <="001011001000"; -- Argumento 2511 Funcion -0.65201053
  when "100111010000"=> s <="001011000110"; -- Argumento 2512 Funcion -0.65317284
  when "100111010001"=> s <="001011000011"; -- Argumento 2513 Funcion -0.65433362
  when "100111010010"=> s <="001011000001"; -- Argumento 2514 Funcion -0.65549285
  when "100111010011"=> s <="001010111111"; -- Argumento 2515 Funcion -0.65665055
  when "100111010100"=> s <="001010111100"; -- Argumento 2516 Funcion -0.65780669
  when "100111010101"=> s <="001010111010"; -- Argumento 2517 Funcion -0.65896129
  when "100111010110"=> s <="001010111000"; -- Argumento 2518 Funcion -0.66011434
  when "100111010111"=> s <="001010110101"; -- Argumento 2519 Funcion -0.66126584
  when "100111011000"=> s <="001010110011"; -- Argumento 2520 Funcion -0.66241578
  when "100111011001"=> s <="001010110001"; -- Argumento 2521 Funcion -0.66356416
  when "100111011010"=> s <="001010101110"; -- Argumento 2522 Funcion -0.66471098
  when "100111011011"=> s <="001010101100"; -- Argumento 2523 Funcion -0.66585623
  when "100111011100"=> s <="001010101001"; -- Argumento 2524 Funcion -0.66699992
  when "100111011101"=> s <="001010100111"; -- Argumento 2525 Funcion -0.66814204
  when "100111011110"=> s <="001010100101"; -- Argumento 2526 Funcion -0.66928259
  when "100111011111"=> s <="001010100010"; -- Argumento 2527 Funcion -0.67042156
  when "100111100000"=> s <="001010100000"; -- Argumento 2528 Funcion -0.67155895
  when "100111100001"=> s <="001010011110"; -- Argumento 2529 Funcion -0.67269477
  when "100111100010"=> s <="001010011011"; -- Argumento 2530 Funcion -0.67382900
  when "100111100011"=> s <="001010011001"; -- Argumento 2531 Funcion -0.67496165
  when "100111100100"=> s <="001010010111"; -- Argumento 2532 Funcion -0.67609270
  when "100111100101"=> s <="001010010101"; -- Argumento 2533 Funcion -0.67722217
  when "100111100110"=> s <="001010010010"; -- Argumento 2534 Funcion -0.67835004
  when "100111100111"=> s <="001010010000"; -- Argumento 2535 Funcion -0.67947632
  when "100111101000"=> s <="001010001110"; -- Argumento 2536 Funcion -0.68060100
  when "100111101001"=> s <="001010001011"; -- Argumento 2537 Funcion -0.68172407
  when "100111101010"=> s <="001010001001"; -- Argumento 2538 Funcion -0.68284555
  when "100111101011"=> s <="001010000111"; -- Argumento 2539 Funcion -0.68396541
  when "100111101100"=> s <="001010000100"; -- Argumento 2540 Funcion -0.68508367
  when "100111101101"=> s <="001010000010"; -- Argumento 2541 Funcion -0.68620031
  when "100111101110"=> s <="001010000000"; -- Argumento 2542 Funcion -0.68731534
  when "100111101111"=> s <="001001111110"; -- Argumento 2543 Funcion -0.68842875
  when "100111110000"=> s <="001001111011"; -- Argumento 2544 Funcion -0.68954054
  when "100111110001"=> s <="001001111001"; -- Argumento 2545 Funcion -0.69065071
  when "100111110010"=> s <="001001110111"; -- Argumento 2546 Funcion -0.69175926
  when "100111110011"=> s <="001001110101"; -- Argumento 2547 Funcion -0.69286617
  when "100111110100"=> s <="001001110010"; -- Argumento 2548 Funcion -0.69397146
  when "100111110101"=> s <="001001110000"; -- Argumento 2549 Funcion -0.69507511
  when "100111110110"=> s <="001001101110"; -- Argumento 2550 Funcion -0.69617713
  when "100111110111"=> s <="001001101011"; -- Argumento 2551 Funcion -0.69727751
  when "100111111000"=> s <="001001101001"; -- Argumento 2552 Funcion -0.69837625
  when "100111111001"=> s <="001001100111"; -- Argumento 2553 Funcion -0.69947334
  when "100111111010"=> s <="001001100101"; -- Argumento 2554 Funcion -0.70056879
  when "100111111011"=> s <="001001100010"; -- Argumento 2555 Funcion -0.70166259
  when "100111111100"=> s <="001001100000"; -- Argumento 2556 Funcion -0.70275474
  when "100111111101"=> s <="001001011110"; -- Argumento 2557 Funcion -0.70384524
  when "100111111110"=> s <="001001011100"; -- Argumento 2558 Funcion -0.70493408
  when "100111111111"=> s <="001001011010"; -- Argumento 2559 Funcion -0.70602126
  when "101000000000"=> s <="001001010111"; -- Argumento 2560 Funcion -0.70710678
  when "101000000001"=> s <="001001010101"; -- Argumento 2561 Funcion -0.70819064
  when "101000000010"=> s <="001001010011"; -- Argumento 2562 Funcion -0.70927283
  when "101000000011"=> s <="001001010001"; -- Argumento 2563 Funcion -0.71035335
  when "101000000100"=> s <="001001001110"; -- Argumento 2564 Funcion -0.71143220
  when "101000000101"=> s <="001001001100"; -- Argumento 2565 Funcion -0.71250937
  when "101000000110"=> s <="001001001010"; -- Argumento 2566 Funcion -0.71358487
  when "101000000111"=> s <="001001001000"; -- Argumento 2567 Funcion -0.71465869
  when "101000001000"=> s <="001001000110"; -- Argumento 2568 Funcion -0.71573083
  when "101000001001"=> s <="001001000011"; -- Argumento 2569 Funcion -0.71680128
  when "101000001010"=> s <="001001000001"; -- Argumento 2570 Funcion -0.71787005
  when "101000001011"=> s <="001000111111"; -- Argumento 2571 Funcion -0.71893712
  when "101000001100"=> s <="001000111101"; -- Argumento 2572 Funcion -0.72000251
  when "101000001101"=> s <="001000111011"; -- Argumento 2573 Funcion -0.72106620
  when "101000001110"=> s <="001000111001"; -- Argumento 2574 Funcion -0.72212819
  when "101000001111"=> s <="001000110110"; -- Argumento 2575 Funcion -0.72318849
  when "101000010000"=> s <="001000110100"; -- Argumento 2576 Funcion -0.72424708
  when "101000010001"=> s <="001000110010"; -- Argumento 2577 Funcion -0.72530397
  when "101000010010"=> s <="001000110000"; -- Argumento 2578 Funcion -0.72635916
  when "101000010011"=> s <="001000101110"; -- Argumento 2579 Funcion -0.72741263
  when "101000010100"=> s <="001000101100"; -- Argumento 2580 Funcion -0.72846439
  when "101000010101"=> s <="001000101001"; -- Argumento 2581 Funcion -0.72951444
  when "101000010110"=> s <="001000100111"; -- Argumento 2582 Funcion -0.73056277
  when "101000010111"=> s <="001000100101"; -- Argumento 2583 Funcion -0.73160938
  when "101000011000"=> s <="001000100011"; -- Argumento 2584 Funcion -0.73265427
  when "101000011001"=> s <="001000100001"; -- Argumento 2585 Funcion -0.73369744
  when "101000011010"=> s <="001000011111"; -- Argumento 2586 Funcion -0.73473888
  when "101000011011"=> s <="001000011101"; -- Argumento 2587 Funcion -0.73577859
  when "101000011100"=> s <="001000011010"; -- Argumento 2588 Funcion -0.73681657
  when "101000011101"=> s <="001000011000"; -- Argumento 2589 Funcion -0.73785281
  when "101000011110"=> s <="001000010110"; -- Argumento 2590 Funcion -0.73888732
  when "101000011111"=> s <="001000010100"; -- Argumento 2591 Funcion -0.73992010
  when "101000100000"=> s <="001000010010"; -- Argumento 2592 Funcion -0.74095113
  when "101000100001"=> s <="001000010000"; -- Argumento 2593 Funcion -0.74198041
  when "101000100010"=> s <="001000001110"; -- Argumento 2594 Funcion -0.74300795
  when "101000100011"=> s <="001000001100"; -- Argumento 2595 Funcion -0.74403374
  when "101000100100"=> s <="001000001010"; -- Argumento 2596 Funcion -0.74505779
  when "101000100101"=> s <="001000001000"; -- Argumento 2597 Funcion -0.74608007
  when "101000100110"=> s <="001000000101"; -- Argumento 2598 Funcion -0.74710061
  when "101000100111"=> s <="001000000011"; -- Argumento 2599 Funcion -0.74811938
  when "101000101000"=> s <="001000000001"; -- Argumento 2600 Funcion -0.74913639
  when "101000101001"=> s <="000111111111"; -- Argumento 2601 Funcion -0.75015165
  when "101000101010"=> s <="000111111101"; -- Argumento 2602 Funcion -0.75116513
  when "101000101011"=> s <="000111111011"; -- Argumento 2603 Funcion -0.75217685
  when "101000101100"=> s <="000111111001"; -- Argumento 2604 Funcion -0.75318680
  when "101000101101"=> s <="000111110111"; -- Argumento 2605 Funcion -0.75419498
  when "101000101110"=> s <="000111110101"; -- Argumento 2606 Funcion -0.75520138
  when "101000101111"=> s <="000111110011"; -- Argumento 2607 Funcion -0.75620600
  when "101000110000"=> s <="000111110001"; -- Argumento 2608 Funcion -0.75720885
  when "101000110001"=> s <="000111101111"; -- Argumento 2609 Funcion -0.75820991
  when "101000110010"=> s <="000111101101"; -- Argumento 2610 Funcion -0.75920919
  when "101000110011"=> s <="000111101011"; -- Argumento 2611 Funcion -0.76020668
  when "101000110100"=> s <="000111101001"; -- Argumento 2612 Funcion -0.76120239
  when "101000110101"=> s <="000111100111"; -- Argumento 2613 Funcion -0.76219630
  when "101000110110"=> s <="000111100100"; -- Argumento 2614 Funcion -0.76318842
  when "101000110111"=> s <="000111100010"; -- Argumento 2615 Funcion -0.76417874
  when "101000111000"=> s <="000111100000"; -- Argumento 2616 Funcion -0.76516727
  when "101000111001"=> s <="000111011110"; -- Argumento 2617 Funcion -0.76615399
  when "101000111010"=> s <="000111011100"; -- Argumento 2618 Funcion -0.76713891
  when "101000111011"=> s <="000111011010"; -- Argumento 2619 Funcion -0.76812203
  when "101000111100"=> s <="000111011000"; -- Argumento 2620 Funcion -0.76910334
  when "101000111101"=> s <="000111010110"; -- Argumento 2621 Funcion -0.77008284
  when "101000111110"=> s <="000111010100"; -- Argumento 2622 Funcion -0.77106052
  when "101000111111"=> s <="000111010010"; -- Argumento 2623 Funcion -0.77203640
  when "101001000000"=> s <="000111010000"; -- Argumento 2624 Funcion -0.77301045
  when "101001000001"=> s <="000111001110"; -- Argumento 2625 Funcion -0.77398269
  when "101001000010"=> s <="000111001100"; -- Argumento 2626 Funcion -0.77495311
  when "101001000011"=> s <="000111001010"; -- Argumento 2627 Funcion -0.77592170
  when "101001000100"=> s <="000111001000"; -- Argumento 2628 Funcion -0.77688847
  when "101001000101"=> s <="000111000110"; -- Argumento 2629 Funcion -0.77785340
  when "101001000110"=> s <="000111000100"; -- Argumento 2630 Funcion -0.77881651
  when "101001000111"=> s <="000111000011"; -- Argumento 2631 Funcion -0.77977779
  when "101001001000"=> s <="000111000001"; -- Argumento 2632 Funcion -0.78073723
  when "101001001001"=> s <="000110111111"; -- Argumento 2633 Funcion -0.78169483
  when "101001001010"=> s <="000110111101"; -- Argumento 2634 Funcion -0.78265060
  when "101001001011"=> s <="000110111011"; -- Argumento 2635 Funcion -0.78360452
  when "101001001100"=> s <="000110111001"; -- Argumento 2636 Funcion -0.78455660
  when "101001001101"=> s <="000110110111"; -- Argumento 2637 Funcion -0.78550683
  when "101001001110"=> s <="000110110101"; -- Argumento 2638 Funcion -0.78645521
  when "101001001111"=> s <="000110110011"; -- Argumento 2639 Funcion -0.78740175
  when "101001010000"=> s <="000110110001"; -- Argumento 2640 Funcion -0.78834643
  when "101001010001"=> s <="000110101111"; -- Argumento 2641 Funcion -0.78928925
  when "101001010010"=> s <="000110101101"; -- Argumento 2642 Funcion -0.79023022
  when "101001010011"=> s <="000110101011"; -- Argumento 2643 Funcion -0.79116933
  when "101001010100"=> s <="000110101001"; -- Argumento 2644 Funcion -0.79210658
  when "101001010101"=> s <="000110100111"; -- Argumento 2645 Funcion -0.79304196
  when "101001010110"=> s <="000110100101"; -- Argumento 2646 Funcion -0.79397548
  when "101001010111"=> s <="000110100100"; -- Argumento 2647 Funcion -0.79490713
  when "101001011000"=> s <="000110100010"; -- Argumento 2648 Funcion -0.79583690
  when "101001011001"=> s <="000110100000"; -- Argumento 2649 Funcion -0.79676481
  when "101001011010"=> s <="000110011110"; -- Argumento 2650 Funcion -0.79769084
  when "101001011011"=> s <="000110011100"; -- Argumento 2651 Funcion -0.79861499
  when "101001011100"=> s <="000110011010"; -- Argumento 2652 Funcion -0.79953727
  when "101001011101"=> s <="000110011000"; -- Argumento 2653 Funcion -0.80045766
  when "101001011110"=> s <="000110010110"; -- Argumento 2654 Funcion -0.80137617
  when "101001011111"=> s <="000110010100"; -- Argumento 2655 Funcion -0.80229280
  when "101001100000"=> s <="000110010011"; -- Argumento 2656 Funcion -0.80320753
  when "101001100001"=> s <="000110010001"; -- Argumento 2657 Funcion -0.80412038
  when "101001100010"=> s <="000110001111"; -- Argumento 2658 Funcion -0.80503133
  when "101001100011"=> s <="000110001101"; -- Argumento 2659 Funcion -0.80594039
  when "101001100100"=> s <="000110001011"; -- Argumento 2660 Funcion -0.80684755
  when "101001100101"=> s <="000110001001"; -- Argumento 2661 Funcion -0.80775282
  when "101001100110"=> s <="000110000111"; -- Argumento 2662 Funcion -0.80865618
  when "101001100111"=> s <="000110000110"; -- Argumento 2663 Funcion -0.80955764
  when "101001101000"=> s <="000110000100"; -- Argumento 2664 Funcion -0.81045720
  when "101001101001"=> s <="000110000010"; -- Argumento 2665 Funcion -0.81135485
  when "101001101010"=> s <="000110000000"; -- Argumento 2666 Funcion -0.81225059
  when "101001101011"=> s <="000101111110"; -- Argumento 2667 Funcion -0.81314441
  when "101001101100"=> s <="000101111100"; -- Argumento 2668 Funcion -0.81403633
  when "101001101101"=> s <="000101111011"; -- Argumento 2669 Funcion -0.81492633
  when "101001101110"=> s <="000101111001"; -- Argumento 2670 Funcion -0.81581441
  when "101001101111"=> s <="000101110111"; -- Argumento 2671 Funcion -0.81670057
  when "101001110000"=> s <="000101110101"; -- Argumento 2672 Funcion -0.81758481
  when "101001110001"=> s <="000101110011"; -- Argumento 2673 Funcion -0.81846713
  when "101001110010"=> s <="000101110001"; -- Argumento 2674 Funcion -0.81934752
  when "101001110011"=> s <="000101110000"; -- Argumento 2675 Funcion -0.82022598
  when "101001110100"=> s <="000101101110"; -- Argumento 2676 Funcion -0.82110251
  when "101001110101"=> s <="000101101100"; -- Argumento 2677 Funcion -0.82197712
  when "101001110110"=> s <="000101101010"; -- Argumento 2678 Funcion -0.82284978
  when "101001110111"=> s <="000101101001"; -- Argumento 2679 Funcion -0.82372051
  when "101001111000"=> s <="000101100111"; -- Argumento 2680 Funcion -0.82458930
  when "101001111001"=> s <="000101100101"; -- Argumento 2681 Funcion -0.82545615
  when "101001111010"=> s <="000101100011"; -- Argumento 2682 Funcion -0.82632106
  when "101001111011"=> s <="000101100001"; -- Argumento 2683 Funcion -0.82718403
  when "101001111100"=> s <="000101100000"; -- Argumento 2684 Funcion -0.82804505
  when "101001111101"=> s <="000101011110"; -- Argumento 2685 Funcion -0.82890411
  when "101001111110"=> s <="000101011100"; -- Argumento 2686 Funcion -0.82976123
  when "101001111111"=> s <="000101011010"; -- Argumento 2687 Funcion -0.83061640
  when "101010000000"=> s <="000101011001"; -- Argumento 2688 Funcion -0.83146961
  when "101010000001"=> s <="000101010111"; -- Argumento 2689 Funcion -0.83232087
  when "101010000010"=> s <="000101010101"; -- Argumento 2690 Funcion -0.83317016
  when "101010000011"=> s <="000101010011"; -- Argumento 2691 Funcion -0.83401750
  when "101010000100"=> s <="000101010010"; -- Argumento 2692 Funcion -0.83486287
  when "101010000101"=> s <="000101010000"; -- Argumento 2693 Funcion -0.83570628
  when "101010000110"=> s <="000101001110"; -- Argumento 2694 Funcion -0.83654773
  when "101010000111"=> s <="000101001101"; -- Argumento 2695 Funcion -0.83738720
  when "101010001000"=> s <="000101001011"; -- Argumento 2696 Funcion -0.83822471
  when "101010001001"=> s <="000101001001"; -- Argumento 2697 Funcion -0.83906024
  when "101010001010"=> s <="000101000111"; -- Argumento 2698 Funcion -0.83989379
  when "101010001011"=> s <="000101000110"; -- Argumento 2699 Funcion -0.84072537
  when "101010001100"=> s <="000101000100"; -- Argumento 2700 Funcion -0.84155498
  when "101010001101"=> s <="000101000010"; -- Argumento 2701 Funcion -0.84238260
  when "101010001110"=> s <="000101000001"; -- Argumento 2702 Funcion -0.84320824
  when "101010001111"=> s <="000100111111"; -- Argumento 2703 Funcion -0.84403190
  when "101010010000"=> s <="000100111101"; -- Argumento 2704 Funcion -0.84485357
  when "101010010001"=> s <="000100111100"; -- Argumento 2705 Funcion -0.84567325
  when "101010010010"=> s <="000100111010"; -- Argumento 2706 Funcion -0.84649094
  when "101010010011"=> s <="000100111000"; -- Argumento 2707 Funcion -0.84730664
  when "101010010100"=> s <="000100110111"; -- Argumento 2708 Funcion -0.84812034
  when "101010010101"=> s <="000100110101"; -- Argumento 2709 Funcion -0.84893206
  when "101010010110"=> s <="000100110011"; -- Argumento 2710 Funcion -0.84974177
  when "101010010111"=> s <="000100110010"; -- Argumento 2711 Funcion -0.85054948
  when "101010011000"=> s <="000100110000"; -- Argumento 2712 Funcion -0.85135519
  when "101010011001"=> s <="000100101110"; -- Argumento 2713 Funcion -0.85215890
  when "101010011010"=> s <="000100101101"; -- Argumento 2714 Funcion -0.85296060
  when "101010011011"=> s <="000100101011"; -- Argumento 2715 Funcion -0.85376030
  when "101010011100"=> s <="000100101001"; -- Argumento 2716 Funcion -0.85455799
  when "101010011101"=> s <="000100101000"; -- Argumento 2717 Funcion -0.85535366
  when "101010011110"=> s <="000100100110"; -- Argumento 2718 Funcion -0.85614733
  when "101010011111"=> s <="000100100100"; -- Argumento 2719 Funcion -0.85693898
  when "101010100000"=> s <="000100100011"; -- Argumento 2720 Funcion -0.85772861
  when "101010100001"=> s <="000100100001"; -- Argumento 2721 Funcion -0.85851622
  when "101010100010"=> s <="000100100000"; -- Argumento 2722 Funcion -0.85930182
  when "101010100011"=> s <="000100011110"; -- Argumento 2723 Funcion -0.86008539
  when "101010100100"=> s <="000100011100"; -- Argumento 2724 Funcion -0.86086694
  when "101010100101"=> s <="000100011011"; -- Argumento 2725 Funcion -0.86164646
  when "101010100110"=> s <="000100011001"; -- Argumento 2726 Funcion -0.86242396
  when "101010100111"=> s <="000100011000"; -- Argumento 2727 Funcion -0.86319942
  when "101010101000"=> s <="000100010110"; -- Argumento 2728 Funcion -0.86397286
  when "101010101001"=> s <="000100010101"; -- Argumento 2729 Funcion -0.86474426
  when "101010101010"=> s <="000100010011"; -- Argumento 2730 Funcion -0.86551362
  when "101010101011"=> s <="000100010001"; -- Argumento 2731 Funcion -0.86628095
  when "101010101100"=> s <="000100010000"; -- Argumento 2732 Funcion -0.86704625
  when "101010101101"=> s <="000100001110"; -- Argumento 2733 Funcion -0.86780950
  when "101010101110"=> s <="000100001101"; -- Argumento 2734 Funcion -0.86857071
  when "101010101111"=> s <="000100001011"; -- Argumento 2735 Funcion -0.86932987
  when "101010110000"=> s <="000100001010"; -- Argumento 2736 Funcion -0.87008699
  when "101010110001"=> s <="000100001000"; -- Argumento 2737 Funcion -0.87084206
  when "101010110010"=> s <="000100000110"; -- Argumento 2738 Funcion -0.87159509
  when "101010110011"=> s <="000100000101"; -- Argumento 2739 Funcion -0.87234606
  when "101010110100"=> s <="000100000011"; -- Argumento 2740 Funcion -0.87309498
  when "101010110101"=> s <="000100000010"; -- Argumento 2741 Funcion -0.87384184
  when "101010110110"=> s <="000100000000"; -- Argumento 2742 Funcion -0.87458665
  when "101010110111"=> s <="000011111111"; -- Argumento 2743 Funcion -0.87532940
  when "101010111000"=> s <="000011111101"; -- Argumento 2744 Funcion -0.87607009
  when "101010111001"=> s <="000011111100"; -- Argumento 2745 Funcion -0.87680872
  when "101010111010"=> s <="000011111010"; -- Argumento 2746 Funcion -0.87754529
  when "101010111011"=> s <="000011111001"; -- Argumento 2747 Funcion -0.87827979
  when "101010111100"=> s <="000011110111"; -- Argumento 2748 Funcion -0.87901223
  when "101010111101"=> s <="000011110110"; -- Argumento 2749 Funcion -0.87974259
  when "101010111110"=> s <="000011110100"; -- Argumento 2750 Funcion -0.88047089
  when "101010111111"=> s <="000011110011"; -- Argumento 2751 Funcion -0.88119711
  when "101011000000"=> s <="000011110001"; -- Argumento 2752 Funcion -0.88192126
  when "101011000001"=> s <="000011110000"; -- Argumento 2753 Funcion -0.88264334
  when "101011000010"=> s <="000011101110"; -- Argumento 2754 Funcion -0.88336334
  when "101011000011"=> s <="000011101101"; -- Argumento 2755 Funcion -0.88408126
  when "101011000100"=> s <="000011101011"; -- Argumento 2756 Funcion -0.88479710
  when "101011000101"=> s <="000011101010"; -- Argumento 2757 Funcion -0.88551086
  when "101011000110"=> s <="000011101001"; -- Argumento 2758 Funcion -0.88622253
  when "101011000111"=> s <="000011100111"; -- Argumento 2759 Funcion -0.88693212
  when "101011001000"=> s <="000011100110"; -- Argumento 2760 Funcion -0.88763962
  when "101011001001"=> s <="000011100100"; -- Argumento 2761 Funcion -0.88834503
  when "101011001010"=> s <="000011100011"; -- Argumento 2762 Funcion -0.88904836
  when "101011001011"=> s <="000011100001"; -- Argumento 2763 Funcion -0.88974959
  when "101011001100"=> s <="000011100000"; -- Argumento 2764 Funcion -0.89044872
  when "101011001101"=> s <="000011011110"; -- Argumento 2765 Funcion -0.89114576
  when "101011001110"=> s <="000011011101"; -- Argumento 2766 Funcion -0.89184071
  when "101011001111"=> s <="000011011100"; -- Argumento 2767 Funcion -0.89253356
  when "101011010000"=> s <="000011011010"; -- Argumento 2768 Funcion -0.89322430
  when "101011010001"=> s <="000011011001"; -- Argumento 2769 Funcion -0.89391295
  when "101011010010"=> s <="000011010111"; -- Argumento 2770 Funcion -0.89459949
  when "101011010011"=> s <="000011010110"; -- Argumento 2771 Funcion -0.89528392
  when "101011010100"=> s <="000011010101"; -- Argumento 2772 Funcion -0.89596625
  when "101011010101"=> s <="000011010011"; -- Argumento 2773 Funcion -0.89664647
  when "101011010110"=> s <="000011010010"; -- Argumento 2774 Funcion -0.89732458
  when "101011010111"=> s <="000011010000"; -- Argumento 2775 Funcion -0.89800058
  when "101011011000"=> s <="000011001111"; -- Argumento 2776 Funcion -0.89867447
  when "101011011001"=> s <="000011001110"; -- Argumento 2777 Funcion -0.89934624
  when "101011011010"=> s <="000011001100"; -- Argumento 2778 Funcion -0.90001589
  when "101011011011"=> s <="000011001011"; -- Argumento 2779 Funcion -0.90068343
  when "101011011100"=> s <="000011001010"; -- Argumento 2780 Funcion -0.90134885
  when "101011011101"=> s <="000011001000"; -- Argumento 2781 Funcion -0.90201214
  when "101011011110"=> s <="000011000111"; -- Argumento 2782 Funcion -0.90267332
  when "101011011111"=> s <="000011000101"; -- Argumento 2783 Funcion -0.90333237
  when "101011100000"=> s <="000011000100"; -- Argumento 2784 Funcion -0.90398929
  when "101011100001"=> s <="000011000011"; -- Argumento 2785 Funcion -0.90464409
  when "101011100010"=> s <="000011000001"; -- Argumento 2786 Funcion -0.90529676
  when "101011100011"=> s <="000011000000"; -- Argumento 2787 Funcion -0.90594730
  when "101011100100"=> s <="000010111111"; -- Argumento 2788 Funcion -0.90659570
  when "101011100101"=> s <="000010111101"; -- Argumento 2789 Funcion -0.90724198
  when "101011100110"=> s <="000010111100"; -- Argumento 2790 Funcion -0.90788612
  when "101011100111"=> s <="000010111011"; -- Argumento 2791 Funcion -0.90852812
  when "101011101000"=> s <="000010111010"; -- Argumento 2792 Funcion -0.90916798
  when "101011101001"=> s <="000010111000"; -- Argumento 2793 Funcion -0.90980571
  when "101011101010"=> s <="000010110111"; -- Argumento 2794 Funcion -0.91044129
  when "101011101011"=> s <="000010110110"; -- Argumento 2795 Funcion -0.91107473
  when "101011101100"=> s <="000010110100"; -- Argumento 2796 Funcion -0.91170603
  when "101011101101"=> s <="000010110011"; -- Argumento 2797 Funcion -0.91233518
  when "101011101110"=> s <="000010110010"; -- Argumento 2798 Funcion -0.91296219
  when "101011101111"=> s <="000010110000"; -- Argumento 2799 Funcion -0.91358705
  when "101011110000"=> s <="000010101111"; -- Argumento 2800 Funcion -0.91420976
  when "101011110001"=> s <="000010101110"; -- Argumento 2801 Funcion -0.91483031
  when "101011110010"=> s <="000010101101"; -- Argumento 2802 Funcion -0.91544872
  when "101011110011"=> s <="000010101011"; -- Argumento 2803 Funcion -0.91606497
  when "101011110100"=> s <="000010101010"; -- Argumento 2804 Funcion -0.91667906
  when "101011110101"=> s <="000010101001"; -- Argumento 2805 Funcion -0.91729100
  when "101011110110"=> s <="000010101000"; -- Argumento 2806 Funcion -0.91790078
  when "101011110111"=> s <="000010100110"; -- Argumento 2807 Funcion -0.91850839
  when "101011111000"=> s <="000010100101"; -- Argumento 2808 Funcion -0.91911385
  when "101011111001"=> s <="000010100100"; -- Argumento 2809 Funcion -0.91971715
  when "101011111010"=> s <="000010100011"; -- Argumento 2810 Funcion -0.92031828
  when "101011111011"=> s <="000010100001"; -- Argumento 2811 Funcion -0.92091724
  when "101011111100"=> s <="000010100000"; -- Argumento 2812 Funcion -0.92151404
  when "101011111101"=> s <="000010011111"; -- Argumento 2813 Funcion -0.92210867
  when "101011111110"=> s <="000010011110"; -- Argumento 2814 Funcion -0.92270113
  when "101011111111"=> s <="000010011101"; -- Argumento 2815 Funcion -0.92329142
  when "101100000000"=> s <="000010011011"; -- Argumento 2816 Funcion -0.92387953
  when "101100000001"=> s <="000010011010"; -- Argumento 2817 Funcion -0.92446547
  when "101100000010"=> s <="000010011001"; -- Argumento 2818 Funcion -0.92504924
  when "101100000011"=> s <="000010011000"; -- Argumento 2819 Funcion -0.92563083
  when "101100000100"=> s <="000010010111"; -- Argumento 2820 Funcion -0.92621024
  when "101100000101"=> s <="000010010101"; -- Argumento 2821 Funcion -0.92678747
  when "101100000110"=> s <="000010010100"; -- Argumento 2822 Funcion -0.92736253
  when "101100000111"=> s <="000010010011"; -- Argumento 2823 Funcion -0.92793539
  when "101100001000"=> s <="000010010010"; -- Argumento 2824 Funcion -0.92850608
  when "101100001001"=> s <="000010010001"; -- Argumento 2825 Funcion -0.92907458
  when "101100001010"=> s <="000010010000"; -- Argumento 2826 Funcion -0.92964090
  when "101100001011"=> s <="000010001110"; -- Argumento 2827 Funcion -0.93020502
  when "101100001100"=> s <="000010001101"; -- Argumento 2828 Funcion -0.93076696
  when "101100001101"=> s <="000010001100"; -- Argumento 2829 Funcion -0.93132671
  when "101100001110"=> s <="000010001011"; -- Argumento 2830 Funcion -0.93188427
  when "101100001111"=> s <="000010001010"; -- Argumento 2831 Funcion -0.93243963
  when "101100010000"=> s <="000010001001"; -- Argumento 2832 Funcion -0.93299280
  when "101100010001"=> s <="000010001000"; -- Argumento 2833 Funcion -0.93354377
  when "101100010010"=> s <="000010000110"; -- Argumento 2834 Funcion -0.93409255
  when "101100010011"=> s <="000010000101"; -- Argumento 2835 Funcion -0.93463913
  when "101100010100"=> s <="000010000100"; -- Argumento 2836 Funcion -0.93518351
  when "101100010101"=> s <="000010000011"; -- Argumento 2837 Funcion -0.93572569
  when "101100010110"=> s <="000010000010"; -- Argumento 2838 Funcion -0.93626567
  when "101100010111"=> s <="000010000001"; -- Argumento 2839 Funcion -0.93680344
  when "101100011000"=> s <="000010000000"; -- Argumento 2840 Funcion -0.93733901
  when "101100011001"=> s <="000001111111"; -- Argumento 2841 Funcion -0.93787238
  when "101100011010"=> s <="000001111110"; -- Argumento 2842 Funcion -0.93840353
  when "101100011011"=> s <="000001111101"; -- Argumento 2843 Funcion -0.93893248
  when "101100011100"=> s <="000001111011"; -- Argumento 2844 Funcion -0.93945922
  when "101100011101"=> s <="000001111010"; -- Argumento 2845 Funcion -0.93998375
  when "101100011110"=> s <="000001111001"; -- Argumento 2846 Funcion -0.94050607
  when "101100011111"=> s <="000001111000"; -- Argumento 2847 Funcion -0.94102618
  when "101100100000"=> s <="000001110111"; -- Argumento 2848 Funcion -0.94154407
  when "101100100001"=> s <="000001110110"; -- Argumento 2849 Funcion -0.94205974
  when "101100100010"=> s <="000001110101"; -- Argumento 2850 Funcion -0.94257320
  when "101100100011"=> s <="000001110100"; -- Argumento 2851 Funcion -0.94308444
  when "101100100100"=> s <="000001110011"; -- Argumento 2852 Funcion -0.94359346
  when "101100100101"=> s <="000001110010"; -- Argumento 2853 Funcion -0.94410026
  when "101100100110"=> s <="000001110001"; -- Argumento 2854 Funcion -0.94460484
  when "101100100111"=> s <="000001110000"; -- Argumento 2855 Funcion -0.94510719
  when "101100101000"=> s <="000001101111"; -- Argumento 2856 Funcion -0.94560733
  when "101100101001"=> s <="000001101110"; -- Argumento 2857 Funcion -0.94610523
  when "101100101010"=> s <="000001101101"; -- Argumento 2858 Funcion -0.94660091
  when "101100101011"=> s <="000001101100"; -- Argumento 2859 Funcion -0.94709437
  when "101100101100"=> s <="000001101011"; -- Argumento 2860 Funcion -0.94758559
  when "101100101101"=> s <="000001101010"; -- Argumento 2861 Funcion -0.94807459
  when "101100101110"=> s <="000001101001"; -- Argumento 2862 Funcion -0.94856135
  when "101100101111"=> s <="000001101000"; -- Argumento 2863 Funcion -0.94904588
  when "101100110000"=> s <="000001100111"; -- Argumento 2864 Funcion -0.94952818
  when "101100110001"=> s <="000001100110"; -- Argumento 2865 Funcion -0.95000825
  when "101100110010"=> s <="000001100101"; -- Argumento 2866 Funcion -0.95048607
  when "101100110011"=> s <="000001100100"; -- Argumento 2867 Funcion -0.95096167
  when "101100110100"=> s <="000001100011"; -- Argumento 2868 Funcion -0.95143502
  when "101100110101"=> s <="000001100010"; -- Argumento 2869 Funcion -0.95190614
  when "101100110110"=> s <="000001100001"; -- Argumento 2870 Funcion -0.95237501
  when "101100110111"=> s <="000001100000"; -- Argumento 2871 Funcion -0.95284165
  when "101100111000"=> s <="000001011111"; -- Argumento 2872 Funcion -0.95330604
  when "101100111001"=> s <="000001011110"; -- Argumento 2873 Funcion -0.95376819
  when "101100111010"=> s <="000001011101"; -- Argumento 2874 Funcion -0.95422810
  when "101100111011"=> s <="000001011100"; -- Argumento 2875 Funcion -0.95468575
  when "101100111100"=> s <="000001011011"; -- Argumento 2876 Funcion -0.95514117
  when "101100111101"=> s <="000001011010"; -- Argumento 2877 Funcion -0.95559433
  when "101100111110"=> s <="000001011010"; -- Argumento 2878 Funcion -0.95604525
  when "101100111111"=> s <="000001011001"; -- Argumento 2879 Funcion -0.95649392
  when "101101000000"=> s <="000001011000"; -- Argumento 2880 Funcion -0.95694034
  when "101101000001"=> s <="000001010111"; -- Argumento 2881 Funcion -0.95738450
  when "101101000010"=> s <="000001010110"; -- Argumento 2882 Funcion -0.95782641
  when "101101000011"=> s <="000001010101"; -- Argumento 2883 Funcion -0.95826607
  when "101101000100"=> s <="000001010100"; -- Argumento 2884 Funcion -0.95870347
  when "101101000101"=> s <="000001010011"; -- Argumento 2885 Funcion -0.95913862
  when "101101000110"=> s <="000001010010"; -- Argumento 2886 Funcion -0.95957151
  when "101101000111"=> s <="000001010001"; -- Argumento 2887 Funcion -0.96000215
  when "101101001000"=> s <="000001010001"; -- Argumento 2888 Funcion -0.96043052
  when "101101001001"=> s <="000001010000"; -- Argumento 2889 Funcion -0.96085663
  when "101101001010"=> s <="000001001111"; -- Argumento 2890 Funcion -0.96128049
  when "101101001011"=> s <="000001001110"; -- Argumento 2891 Funcion -0.96170208
  when "101101001100"=> s <="000001001101"; -- Argumento 2892 Funcion -0.96212140
  when "101101001101"=> s <="000001001100"; -- Argumento 2893 Funcion -0.96253847
  when "101101001110"=> s <="000001001011"; -- Argumento 2894 Funcion -0.96295327
  when "101101001111"=> s <="000001001011"; -- Argumento 2895 Funcion -0.96336580
  when "101101010000"=> s <="000001001010"; -- Argumento 2896 Funcion -0.96377607
  when "101101010001"=> s <="000001001001"; -- Argumento 2897 Funcion -0.96418406
  when "101101010010"=> s <="000001001000"; -- Argumento 2898 Funcion -0.96458979
  when "101101010011"=> s <="000001000111"; -- Argumento 2899 Funcion -0.96499325
  when "101101010100"=> s <="000001000110"; -- Argumento 2900 Funcion -0.96539444
  when "101101010101"=> s <="000001000110"; -- Argumento 2901 Funcion -0.96579336
  when "101101010110"=> s <="000001000101"; -- Argumento 2902 Funcion -0.96619000
  when "101101010111"=> s <="000001000100"; -- Argumento 2903 Funcion -0.96658437
  when "101101011000"=> s <="000001000011"; -- Argumento 2904 Funcion -0.96697647
  when "101101011001"=> s <="000001000010"; -- Argumento 2905 Funcion -0.96736629
  when "101101011010"=> s <="000001000010"; -- Argumento 2906 Funcion -0.96775384
  when "101101011011"=> s <="000001000001"; -- Argumento 2907 Funcion -0.96813910
  when "101101011100"=> s <="000001000000"; -- Argumento 2908 Funcion -0.96852209
  when "101101011101"=> s <="000000111111"; -- Argumento 2909 Funcion -0.96890280
  when "101101011110"=> s <="000000111110"; -- Argumento 2910 Funcion -0.96928124
  when "101101011111"=> s <="000000111110"; -- Argumento 2911 Funcion -0.96965739
  when "101101100000"=> s <="000000111101"; -- Argumento 2912 Funcion -0.97003125
  when "101101100001"=> s <="000000111100"; -- Argumento 2913 Funcion -0.97040284
  when "101101100010"=> s <="000000111011"; -- Argumento 2914 Funcion -0.97077214
  when "101101100011"=> s <="000000111011"; -- Argumento 2915 Funcion -0.97113916
  when "101101100100"=> s <="000000111010"; -- Argumento 2916 Funcion -0.97150389
  when "101101100101"=> s <="000000111001"; -- Argumento 2917 Funcion -0.97186634
  when "101101100110"=> s <="000000111000"; -- Argumento 2918 Funcion -0.97222650
  when "101101100111"=> s <="000000111000"; -- Argumento 2919 Funcion -0.97258437
  when "101101101000"=> s <="000000110111"; -- Argumento 2920 Funcion -0.97293995
  when "101101101001"=> s <="000000110110"; -- Argumento 2921 Funcion -0.97329325
  when "101101101010"=> s <="000000110101"; -- Argumento 2922 Funcion -0.97364425
  when "101101101011"=> s <="000000110101"; -- Argumento 2923 Funcion -0.97399296
  when "101101101100"=> s <="000000110100"; -- Argumento 2924 Funcion -0.97433938
  when "101101101101"=> s <="000000110011"; -- Argumento 2925 Funcion -0.97468351
  when "101101101110"=> s <="000000110011"; -- Argumento 2926 Funcion -0.97502535
  when "101101101111"=> s <="000000110010"; -- Argumento 2927 Funcion -0.97536489
  when "101101110000"=> s <="000000110001"; -- Argumento 2928 Funcion -0.97570213
  when "101101110001"=> s <="000000110001"; -- Argumento 2929 Funcion -0.97603708
  when "101101110010"=> s <="000000110000"; -- Argumento 2930 Funcion -0.97636973
  when "101101110011"=> s <="000000101111"; -- Argumento 2931 Funcion -0.97670009
  when "101101110100"=> s <="000000101111"; -- Argumento 2932 Funcion -0.97702814
  when "101101110101"=> s <="000000101110"; -- Argumento 2933 Funcion -0.97735390
  when "101101110110"=> s <="000000101101"; -- Argumento 2934 Funcion -0.97767736
  when "101101110111"=> s <="000000101101"; -- Argumento 2935 Funcion -0.97799851
  when "101101111000"=> s <="000000101100"; -- Argumento 2936 Funcion -0.97831737
  when "101101111001"=> s <="000000101011"; -- Argumento 2937 Funcion -0.97863392
  when "101101111010"=> s <="000000101011"; -- Argumento 2938 Funcion -0.97894818
  when "101101111011"=> s <="000000101010"; -- Argumento 2939 Funcion -0.97926012
  when "101101111100"=> s <="000000101001"; -- Argumento 2940 Funcion -0.97956977
  when "101101111101"=> s <="000000101001"; -- Argumento 2941 Funcion -0.97987710
  when "101101111110"=> s <="000000101000"; -- Argumento 2942 Funcion -0.98018214
  when "101101111111"=> s <="000000100111"; -- Argumento 2943 Funcion -0.98048486
  when "101110000000"=> s <="000000100111"; -- Argumento 2944 Funcion -0.98078528
  when "101110000001"=> s <="000000100110"; -- Argumento 2945 Funcion -0.98108339
  when "101110000010"=> s <="000000100110"; -- Argumento 2946 Funcion -0.98137919
  when "101110000011"=> s <="000000100101"; -- Argumento 2947 Funcion -0.98167269
  when "101110000100"=> s <="000000100100"; -- Argumento 2948 Funcion -0.98196387
  when "101110000101"=> s <="000000100100"; -- Argumento 2949 Funcion -0.98225274
  when "101110000110"=> s <="000000100011"; -- Argumento 2950 Funcion -0.98253930
  when "101110000111"=> s <="000000100011"; -- Argumento 2951 Funcion -0.98282355
  when "101110001000"=> s <="000000100010"; -- Argumento 2952 Funcion -0.98310549
  when "101110001001"=> s <="000000100010"; -- Argumento 2953 Funcion -0.98338511
  when "101110001010"=> s <="000000100001"; -- Argumento 2954 Funcion -0.98366242
  when "101110001011"=> s <="000000100000"; -- Argumento 2955 Funcion -0.98393741
  when "101110001100"=> s <="000000100000"; -- Argumento 2956 Funcion -0.98421009
  when "101110001101"=> s <="000000011111"; -- Argumento 2957 Funcion -0.98448046
  when "101110001110"=> s <="000000011111"; -- Argumento 2958 Funcion -0.98474850
  when "101110001111"=> s <="000000011110"; -- Argumento 2959 Funcion -0.98501423
  when "101110010000"=> s <="000000011110"; -- Argumento 2960 Funcion -0.98527764
  when "101110010001"=> s <="000000011101"; -- Argumento 2961 Funcion -0.98553874
  when "101110010010"=> s <="000000011101"; -- Argumento 2962 Funcion -0.98579751
  when "101110010011"=> s <="000000011100"; -- Argumento 2963 Funcion -0.98605396
  when "101110010100"=> s <="000000011100"; -- Argumento 2964 Funcion -0.98630810
  when "101110010101"=> s <="000000011011"; -- Argumento 2965 Funcion -0.98655991
  when "101110010110"=> s <="000000011011"; -- Argumento 2966 Funcion -0.98680940
  when "101110010111"=> s <="000000011010"; -- Argumento 2967 Funcion -0.98705657
  when "101110011000"=> s <="000000011010"; -- Argumento 2968 Funcion -0.98730142
  when "101110011001"=> s <="000000011001"; -- Argumento 2969 Funcion -0.98754394
  when "101110011010"=> s <="000000011001"; -- Argumento 2970 Funcion -0.98778414
  when "101110011011"=> s <="000000011000"; -- Argumento 2971 Funcion -0.98802202
  when "101110011100"=> s <="000000011000"; -- Argumento 2972 Funcion -0.98825757
  when "101110011101"=> s <="000000010111"; -- Argumento 2973 Funcion -0.98849079
  when "101110011110"=> s <="000000010111"; -- Argumento 2974 Funcion -0.98872169
  when "101110011111"=> s <="000000010110"; -- Argumento 2975 Funcion -0.98895026
  when "101110100000"=> s <="000000010110"; -- Argumento 2976 Funcion -0.98917651
  when "101110100001"=> s <="000000010101"; -- Argumento 2977 Funcion -0.98940043
  when "101110100010"=> s <="000000010101"; -- Argumento 2978 Funcion -0.98962202
  when "101110100011"=> s <="000000010100"; -- Argumento 2979 Funcion -0.98984128
  when "101110100100"=> s <="000000010100"; -- Argumento 2980 Funcion -0.99005821
  when "101110100101"=> s <="000000010011"; -- Argumento 2981 Funcion -0.99027281
  when "101110100110"=> s <="000000010011"; -- Argumento 2982 Funcion -0.99048508
  when "101110100111"=> s <="000000010011"; -- Argumento 2983 Funcion -0.99069503
  when "101110101000"=> s <="000000010010"; -- Argumento 2984 Funcion -0.99090264
  when "101110101001"=> s <="000000010010"; -- Argumento 2985 Funcion -0.99110791
  when "101110101010"=> s <="000000010001"; -- Argumento 2986 Funcion -0.99131086
  when "101110101011"=> s <="000000010001"; -- Argumento 2987 Funcion -0.99151147
  when "101110101100"=> s <="000000010000"; -- Argumento 2988 Funcion -0.99170975
  when "101110101101"=> s <="000000010000"; -- Argumento 2989 Funcion -0.99190570
  when "101110101110"=> s <="000000010000"; -- Argumento 2990 Funcion -0.99209931
  when "101110101111"=> s <="000000001111"; -- Argumento 2991 Funcion -0.99229059
  when "101110110000"=> s <="000000001111"; -- Argumento 2992 Funcion -0.99247953
  when "101110110001"=> s <="000000001111"; -- Argumento 2993 Funcion -0.99266614
  when "101110110010"=> s <="000000001110"; -- Argumento 2994 Funcion -0.99285041
  when "101110110011"=> s <="000000001110"; -- Argumento 2995 Funcion -0.99303235
  when "101110110100"=> s <="000000001101"; -- Argumento 2996 Funcion -0.99321195
  when "101110110101"=> s <="000000001101"; -- Argumento 2997 Funcion -0.99338921
  when "101110110110"=> s <="000000001101"; -- Argumento 2998 Funcion -0.99356414
  when "101110110111"=> s <="000000001100"; -- Argumento 2999 Funcion -0.99373672
  when "101110111000"=> s <="000000001100"; -- Argumento 3000 Funcion -0.99390697
  when "101110111001"=> s <="000000001100"; -- Argumento 3001 Funcion -0.99407488
  when "101110111010"=> s <="000000001011"; -- Argumento 3002 Funcion -0.99424045
  when "101110111011"=> s <="000000001011"; -- Argumento 3003 Funcion -0.99440368
  when "101110111100"=> s <="000000001011"; -- Argumento 3004 Funcion -0.99456457
  when "101110111101"=> s <="000000001010"; -- Argumento 3005 Funcion -0.99472312
  when "101110111110"=> s <="000000001010"; -- Argumento 3006 Funcion -0.99487933
  when "101110111111"=> s <="000000001010"; -- Argumento 3007 Funcion -0.99503320
  when "101111000000"=> s <="000000001001"; -- Argumento 3008 Funcion -0.99518473
  when "101111000001"=> s <="000000001001"; -- Argumento 3009 Funcion -0.99533391
  when "101111000010"=> s <="000000001001"; -- Argumento 3010 Funcion -0.99548076
  when "101111000011"=> s <="000000001000"; -- Argumento 3011 Funcion -0.99562526
  when "101111000100"=> s <="000000001000"; -- Argumento 3012 Funcion -0.99576741
  when "101111000101"=> s <="000000001000"; -- Argumento 3013 Funcion -0.99590723
  when "101111000110"=> s <="000000001000"; -- Argumento 3014 Funcion -0.99604470
  when "101111000111"=> s <="000000000111"; -- Argumento 3015 Funcion -0.99617983
  when "101111001000"=> s <="000000000111"; -- Argumento 3016 Funcion -0.99631261
  when "101111001001"=> s <="000000000111"; -- Argumento 3017 Funcion -0.99644305
  when "101111001010"=> s <="000000000111"; -- Argumento 3018 Funcion -0.99657115
  when "101111001011"=> s <="000000000110"; -- Argumento 3019 Funcion -0.99669690
  when "101111001100"=> s <="000000000110"; -- Argumento 3020 Funcion -0.99682030
  when "101111001101"=> s <="000000000110"; -- Argumento 3021 Funcion -0.99694136
  when "101111001110"=> s <="000000000110"; -- Argumento 3022 Funcion -0.99706007
  when "101111001111"=> s <="000000000101"; -- Argumento 3023 Funcion -0.99717644
  when "101111010000"=> s <="000000000101"; -- Argumento 3024 Funcion -0.99729046
  when "101111010001"=> s <="000000000101"; -- Argumento 3025 Funcion -0.99740213
  when "101111010010"=> s <="000000000101"; -- Argumento 3026 Funcion -0.99751146
  when "101111010011"=> s <="000000000100"; -- Argumento 3027 Funcion -0.99761844
  when "101111010100"=> s <="000000000100"; -- Argumento 3028 Funcion -0.99772307
  when "101111010101"=> s <="000000000100"; -- Argumento 3029 Funcion -0.99782535
  when "101111010110"=> s <="000000000100"; -- Argumento 3030 Funcion -0.99792529
  when "101111010111"=> s <="000000000100"; -- Argumento 3031 Funcion -0.99802287
  when "101111011000"=> s <="000000000011"; -- Argumento 3032 Funcion -0.99811811
  when "101111011001"=> s <="000000000011"; -- Argumento 3033 Funcion -0.99821100
  when "101111011010"=> s <="000000000011"; -- Argumento 3034 Funcion -0.99830154
  when "101111011011"=> s <="000000000011"; -- Argumento 3035 Funcion -0.99838974
  when "101111011100"=> s <="000000000011"; -- Argumento 3036 Funcion -0.99847558
  when "101111011101"=> s <="000000000010"; -- Argumento 3037 Funcion -0.99855907
  when "101111011110"=> s <="000000000010"; -- Argumento 3038 Funcion -0.99864022
  when "101111011111"=> s <="000000000010"; -- Argumento 3039 Funcion -0.99871901
  when "101111100000"=> s <="000000000010"; -- Argumento 3040 Funcion -0.99879546
  when "101111100001"=> s <="000000000010"; -- Argumento 3041 Funcion -0.99886955
  when "101111100010"=> s <="000000000010"; -- Argumento 3042 Funcion -0.99894129
  when "101111100011"=> s <="000000000010"; -- Argumento 3043 Funcion -0.99901069
  when "101111100100"=> s <="000000000001"; -- Argumento 3044 Funcion -0.99907773
  when "101111100101"=> s <="000000000001"; -- Argumento 3045 Funcion -0.99914242
  when "101111100110"=> s <="000000000001"; -- Argumento 3046 Funcion -0.99920476
  when "101111100111"=> s <="000000000001"; -- Argumento 3047 Funcion -0.99926475
  when "101111101000"=> s <="000000000001"; -- Argumento 3048 Funcion -0.99932238
  when "101111101001"=> s <="000000000001"; -- Argumento 3049 Funcion -0.99937767
  when "101111101010"=> s <="000000000001"; -- Argumento 3050 Funcion -0.99943060
  when "101111101011"=> s <="000000000001"; -- Argumento 3051 Funcion -0.99948119
  when "101111101100"=> s <="000000000000"; -- Argumento 3052 Funcion -0.99952942
  when "101111101101"=> s <="000000000000"; -- Argumento 3053 Funcion -0.99957530
  when "101111101110"=> s <="000000000000"; -- Argumento 3054 Funcion -0.99961882
  when "101111101111"=> s <="000000000000"; -- Argumento 3055 Funcion -0.99966000
  when "101111110000"=> s <="000000000000"; -- Argumento 3056 Funcion -0.99969882
  when "101111110001"=> s <="000000000000"; -- Argumento 3057 Funcion -0.99973529
  when "101111110010"=> s <="000000000000"; -- Argumento 3058 Funcion -0.99976941
  when "101111110011"=> s <="000000000000"; -- Argumento 3059 Funcion -0.99980117
  when "101111110100"=> s <="000000000000"; -- Argumento 3060 Funcion -0.99983058
  when "101111110101"=> s <="000000000000"; -- Argumento 3061 Funcion -0.99985764
  when "101111110110"=> s <="000000000000"; -- Argumento 3062 Funcion -0.99988235
  when "101111110111"=> s <="000000000000"; -- Argumento 3063 Funcion -0.99990470
  when "101111111000"=> s <="000000000000"; -- Argumento 3064 Funcion -0.99992470
  when "101111111001"=> s <="000000000000"; -- Argumento 3065 Funcion -0.99994235
  when "101111111010"=> s <="000000000000"; -- Argumento 3066 Funcion -0.99995764
  when "101111111011"=> s <="000000000000"; -- Argumento 3067 Funcion -0.99997059
  when "101111111100"=> s <="000000000000"; -- Argumento 3068 Funcion -0.99998118
  when "101111111101"=> s <="000000000000"; -- Argumento 3069 Funcion -0.99998941
  when "101111111110"=> s <="000000000000"; -- Argumento 3070 Funcion -0.99999529
  when "101111111111"=> s <="000000000000"; -- Argumento 3071 Funcion -0.99999882
  when "110000000000"=> s <="000000000000"; -- Argumento 3072 Funcion -1.00000000
  when "110000000001"=> s <="000000000000"; -- Argumento 3073 Funcion -0.99999882
  when "110000000010"=> s <="000000000000"; -- Argumento 3074 Funcion -0.99999529
  when "110000000011"=> s <="000000000000"; -- Argumento 3075 Funcion -0.99998941
  when "110000000100"=> s <="000000000000"; -- Argumento 3076 Funcion -0.99998118
  when "110000000101"=> s <="000000000000"; -- Argumento 3077 Funcion -0.99997059
  when "110000000110"=> s <="000000000000"; -- Argumento 3078 Funcion -0.99995764
  when "110000000111"=> s <="000000000000"; -- Argumento 3079 Funcion -0.99994235
  when "110000001000"=> s <="000000000000"; -- Argumento 3080 Funcion -0.99992470
  when "110000001001"=> s <="000000000000"; -- Argumento 3081 Funcion -0.99990470
  when "110000001010"=> s <="000000000000"; -- Argumento 3082 Funcion -0.99988235
  when "110000001011"=> s <="000000000000"; -- Argumento 3083 Funcion -0.99985764
  when "110000001100"=> s <="000000000000"; -- Argumento 3084 Funcion -0.99983058
  when "110000001101"=> s <="000000000000"; -- Argumento 3085 Funcion -0.99980117
  when "110000001110"=> s <="000000000000"; -- Argumento 3086 Funcion -0.99976941
  when "110000001111"=> s <="000000000000"; -- Argumento 3087 Funcion -0.99973529
  when "110000010000"=> s <="000000000000"; -- Argumento 3088 Funcion -0.99969882
  when "110000010001"=> s <="000000000000"; -- Argumento 3089 Funcion -0.99966000
  when "110000010010"=> s <="000000000000"; -- Argumento 3090 Funcion -0.99961882
  when "110000010011"=> s <="000000000000"; -- Argumento 3091 Funcion -0.99957530
  when "110000010100"=> s <="000000000000"; -- Argumento 3092 Funcion -0.99952942
  when "110000010101"=> s <="000000000001"; -- Argumento 3093 Funcion -0.99948119
  when "110000010110"=> s <="000000000001"; -- Argumento 3094 Funcion -0.99943060
  when "110000010111"=> s <="000000000001"; -- Argumento 3095 Funcion -0.99937767
  when "110000011000"=> s <="000000000001"; -- Argumento 3096 Funcion -0.99932238
  when "110000011001"=> s <="000000000001"; -- Argumento 3097 Funcion -0.99926475
  when "110000011010"=> s <="000000000001"; -- Argumento 3098 Funcion -0.99920476
  when "110000011011"=> s <="000000000001"; -- Argumento 3099 Funcion -0.99914242
  when "110000011100"=> s <="000000000001"; -- Argumento 3100 Funcion -0.99907773
  when "110000011101"=> s <="000000000010"; -- Argumento 3101 Funcion -0.99901069
  when "110000011110"=> s <="000000000010"; -- Argumento 3102 Funcion -0.99894129
  when "110000011111"=> s <="000000000010"; -- Argumento 3103 Funcion -0.99886955
  when "110000100000"=> s <="000000000010"; -- Argumento 3104 Funcion -0.99879546
  when "110000100001"=> s <="000000000010"; -- Argumento 3105 Funcion -0.99871901
  when "110000100010"=> s <="000000000010"; -- Argumento 3106 Funcion -0.99864022
  when "110000100011"=> s <="000000000010"; -- Argumento 3107 Funcion -0.99855907
  when "110000100100"=> s <="000000000011"; -- Argumento 3108 Funcion -0.99847558
  when "110000100101"=> s <="000000000011"; -- Argumento 3109 Funcion -0.99838974
  when "110000100110"=> s <="000000000011"; -- Argumento 3110 Funcion -0.99830154
  when "110000100111"=> s <="000000000011"; -- Argumento 3111 Funcion -0.99821100
  when "110000101000"=> s <="000000000011"; -- Argumento 3112 Funcion -0.99811811
  when "110000101001"=> s <="000000000100"; -- Argumento 3113 Funcion -0.99802287
  when "110000101010"=> s <="000000000100"; -- Argumento 3114 Funcion -0.99792529
  when "110000101011"=> s <="000000000100"; -- Argumento 3115 Funcion -0.99782535
  when "110000101100"=> s <="000000000100"; -- Argumento 3116 Funcion -0.99772307
  when "110000101101"=> s <="000000000100"; -- Argumento 3117 Funcion -0.99761844
  when "110000101110"=> s <="000000000101"; -- Argumento 3118 Funcion -0.99751146
  when "110000101111"=> s <="000000000101"; -- Argumento 3119 Funcion -0.99740213
  when "110000110000"=> s <="000000000101"; -- Argumento 3120 Funcion -0.99729046
  when "110000110001"=> s <="000000000101"; -- Argumento 3121 Funcion -0.99717644
  when "110000110010"=> s <="000000000110"; -- Argumento 3122 Funcion -0.99706007
  when "110000110011"=> s <="000000000110"; -- Argumento 3123 Funcion -0.99694136
  when "110000110100"=> s <="000000000110"; -- Argumento 3124 Funcion -0.99682030
  when "110000110101"=> s <="000000000110"; -- Argumento 3125 Funcion -0.99669690
  when "110000110110"=> s <="000000000111"; -- Argumento 3126 Funcion -0.99657115
  when "110000110111"=> s <="000000000111"; -- Argumento 3127 Funcion -0.99644305
  when "110000111000"=> s <="000000000111"; -- Argumento 3128 Funcion -0.99631261
  when "110000111001"=> s <="000000000111"; -- Argumento 3129 Funcion -0.99617983
  when "110000111010"=> s <="000000001000"; -- Argumento 3130 Funcion -0.99604470
  when "110000111011"=> s <="000000001000"; -- Argumento 3131 Funcion -0.99590723
  when "110000111100"=> s <="000000001000"; -- Argumento 3132 Funcion -0.99576741
  when "110000111101"=> s <="000000001000"; -- Argumento 3133 Funcion -0.99562526
  when "110000111110"=> s <="000000001001"; -- Argumento 3134 Funcion -0.99548076
  when "110000111111"=> s <="000000001001"; -- Argumento 3135 Funcion -0.99533391
  when "110001000000"=> s <="000000001001"; -- Argumento 3136 Funcion -0.99518473
  when "110001000001"=> s <="000000001010"; -- Argumento 3137 Funcion -0.99503320
  when "110001000010"=> s <="000000001010"; -- Argumento 3138 Funcion -0.99487933
  when "110001000011"=> s <="000000001010"; -- Argumento 3139 Funcion -0.99472312
  when "110001000100"=> s <="000000001011"; -- Argumento 3140 Funcion -0.99456457
  when "110001000101"=> s <="000000001011"; -- Argumento 3141 Funcion -0.99440368
  when "110001000110"=> s <="000000001011"; -- Argumento 3142 Funcion -0.99424045
  when "110001000111"=> s <="000000001100"; -- Argumento 3143 Funcion -0.99407488
  when "110001001000"=> s <="000000001100"; -- Argumento 3144 Funcion -0.99390697
  when "110001001001"=> s <="000000001100"; -- Argumento 3145 Funcion -0.99373672
  when "110001001010"=> s <="000000001101"; -- Argumento 3146 Funcion -0.99356414
  when "110001001011"=> s <="000000001101"; -- Argumento 3147 Funcion -0.99338921
  when "110001001100"=> s <="000000001101"; -- Argumento 3148 Funcion -0.99321195
  when "110001001101"=> s <="000000001110"; -- Argumento 3149 Funcion -0.99303235
  when "110001001110"=> s <="000000001110"; -- Argumento 3150 Funcion -0.99285041
  when "110001001111"=> s <="000000001111"; -- Argumento 3151 Funcion -0.99266614
  when "110001010000"=> s <="000000001111"; -- Argumento 3152 Funcion -0.99247953
  when "110001010001"=> s <="000000001111"; -- Argumento 3153 Funcion -0.99229059
  when "110001010010"=> s <="000000010000"; -- Argumento 3154 Funcion -0.99209931
  when "110001010011"=> s <="000000010000"; -- Argumento 3155 Funcion -0.99190570
  when "110001010100"=> s <="000000010000"; -- Argumento 3156 Funcion -0.99170975
  when "110001010101"=> s <="000000010001"; -- Argumento 3157 Funcion -0.99151147
  when "110001010110"=> s <="000000010001"; -- Argumento 3158 Funcion -0.99131086
  when "110001010111"=> s <="000000010010"; -- Argumento 3159 Funcion -0.99110791
  when "110001011000"=> s <="000000010010"; -- Argumento 3160 Funcion -0.99090264
  when "110001011001"=> s <="000000010011"; -- Argumento 3161 Funcion -0.99069503
  when "110001011010"=> s <="000000010011"; -- Argumento 3162 Funcion -0.99048508
  when "110001011011"=> s <="000000010011"; -- Argumento 3163 Funcion -0.99027281
  when "110001011100"=> s <="000000010100"; -- Argumento 3164 Funcion -0.99005821
  when "110001011101"=> s <="000000010100"; -- Argumento 3165 Funcion -0.98984128
  when "110001011110"=> s <="000000010101"; -- Argumento 3166 Funcion -0.98962202
  when "110001011111"=> s <="000000010101"; -- Argumento 3167 Funcion -0.98940043
  when "110001100000"=> s <="000000010110"; -- Argumento 3168 Funcion -0.98917651
  when "110001100001"=> s <="000000010110"; -- Argumento 3169 Funcion -0.98895026
  when "110001100010"=> s <="000000010111"; -- Argumento 3170 Funcion -0.98872169
  when "110001100011"=> s <="000000010111"; -- Argumento 3171 Funcion -0.98849079
  when "110001100100"=> s <="000000011000"; -- Argumento 3172 Funcion -0.98825757
  when "110001100101"=> s <="000000011000"; -- Argumento 3173 Funcion -0.98802202
  when "110001100110"=> s <="000000011001"; -- Argumento 3174 Funcion -0.98778414
  when "110001100111"=> s <="000000011001"; -- Argumento 3175 Funcion -0.98754394
  when "110001101000"=> s <="000000011010"; -- Argumento 3176 Funcion -0.98730142
  when "110001101001"=> s <="000000011010"; -- Argumento 3177 Funcion -0.98705657
  when "110001101010"=> s <="000000011011"; -- Argumento 3178 Funcion -0.98680940
  when "110001101011"=> s <="000000011011"; -- Argumento 3179 Funcion -0.98655991
  when "110001101100"=> s <="000000011100"; -- Argumento 3180 Funcion -0.98630810
  when "110001101101"=> s <="000000011100"; -- Argumento 3181 Funcion -0.98605396
  when "110001101110"=> s <="000000011101"; -- Argumento 3182 Funcion -0.98579751
  when "110001101111"=> s <="000000011101"; -- Argumento 3183 Funcion -0.98553874
  when "110001110000"=> s <="000000011110"; -- Argumento 3184 Funcion -0.98527764
  when "110001110001"=> s <="000000011110"; -- Argumento 3185 Funcion -0.98501423
  when "110001110010"=> s <="000000011111"; -- Argumento 3186 Funcion -0.98474850
  when "110001110011"=> s <="000000011111"; -- Argumento 3187 Funcion -0.98448046
  when "110001110100"=> s <="000000100000"; -- Argumento 3188 Funcion -0.98421009
  when "110001110101"=> s <="000000100000"; -- Argumento 3189 Funcion -0.98393741
  when "110001110110"=> s <="000000100001"; -- Argumento 3190 Funcion -0.98366242
  when "110001110111"=> s <="000000100010"; -- Argumento 3191 Funcion -0.98338511
  when "110001111000"=> s <="000000100010"; -- Argumento 3192 Funcion -0.98310549
  when "110001111001"=> s <="000000100011"; -- Argumento 3193 Funcion -0.98282355
  when "110001111010"=> s <="000000100011"; -- Argumento 3194 Funcion -0.98253930
  when "110001111011"=> s <="000000100100"; -- Argumento 3195 Funcion -0.98225274
  when "110001111100"=> s <="000000100100"; -- Argumento 3196 Funcion -0.98196387
  when "110001111101"=> s <="000000100101"; -- Argumento 3197 Funcion -0.98167269
  when "110001111110"=> s <="000000100110"; -- Argumento 3198 Funcion -0.98137919
  when "110001111111"=> s <="000000100110"; -- Argumento 3199 Funcion -0.98108339
  when "110010000000"=> s <="000000100111"; -- Argumento 3200 Funcion -0.98078528
  when "110010000001"=> s <="000000100111"; -- Argumento 3201 Funcion -0.98048486
  when "110010000010"=> s <="000000101000"; -- Argumento 3202 Funcion -0.98018214
  when "110010000011"=> s <="000000101001"; -- Argumento 3203 Funcion -0.97987710
  when "110010000100"=> s <="000000101001"; -- Argumento 3204 Funcion -0.97956977
  when "110010000101"=> s <="000000101010"; -- Argumento 3205 Funcion -0.97926012
  when "110010000110"=> s <="000000101011"; -- Argumento 3206 Funcion -0.97894818
  when "110010000111"=> s <="000000101011"; -- Argumento 3207 Funcion -0.97863392
  when "110010001000"=> s <="000000101100"; -- Argumento 3208 Funcion -0.97831737
  when "110010001001"=> s <="000000101101"; -- Argumento 3209 Funcion -0.97799851
  when "110010001010"=> s <="000000101101"; -- Argumento 3210 Funcion -0.97767736
  when "110010001011"=> s <="000000101110"; -- Argumento 3211 Funcion -0.97735390
  when "110010001100"=> s <="000000101111"; -- Argumento 3212 Funcion -0.97702814
  when "110010001101"=> s <="000000101111"; -- Argumento 3213 Funcion -0.97670009
  when "110010001110"=> s <="000000110000"; -- Argumento 3214 Funcion -0.97636973
  when "110010001111"=> s <="000000110001"; -- Argumento 3215 Funcion -0.97603708
  when "110010010000"=> s <="000000110001"; -- Argumento 3216 Funcion -0.97570213
  when "110010010001"=> s <="000000110010"; -- Argumento 3217 Funcion -0.97536489
  when "110010010010"=> s <="000000110011"; -- Argumento 3218 Funcion -0.97502535
  when "110010010011"=> s <="000000110011"; -- Argumento 3219 Funcion -0.97468351
  when "110010010100"=> s <="000000110100"; -- Argumento 3220 Funcion -0.97433938
  when "110010010101"=> s <="000000110101"; -- Argumento 3221 Funcion -0.97399296
  when "110010010110"=> s <="000000110101"; -- Argumento 3222 Funcion -0.97364425
  when "110010010111"=> s <="000000110110"; -- Argumento 3223 Funcion -0.97329325
  when "110010011000"=> s <="000000110111"; -- Argumento 3224 Funcion -0.97293995
  when "110010011001"=> s <="000000111000"; -- Argumento 3225 Funcion -0.97258437
  when "110010011010"=> s <="000000111000"; -- Argumento 3226 Funcion -0.97222650
  when "110010011011"=> s <="000000111001"; -- Argumento 3227 Funcion -0.97186634
  when "110010011100"=> s <="000000111010"; -- Argumento 3228 Funcion -0.97150389
  when "110010011101"=> s <="000000111011"; -- Argumento 3229 Funcion -0.97113916
  when "110010011110"=> s <="000000111011"; -- Argumento 3230 Funcion -0.97077214
  when "110010011111"=> s <="000000111100"; -- Argumento 3231 Funcion -0.97040284
  when "110010100000"=> s <="000000111101"; -- Argumento 3232 Funcion -0.97003125
  when "110010100001"=> s <="000000111110"; -- Argumento 3233 Funcion -0.96965739
  when "110010100010"=> s <="000000111110"; -- Argumento 3234 Funcion -0.96928124
  when "110010100011"=> s <="000000111111"; -- Argumento 3235 Funcion -0.96890280
  when "110010100100"=> s <="000001000000"; -- Argumento 3236 Funcion -0.96852209
  when "110010100101"=> s <="000001000001"; -- Argumento 3237 Funcion -0.96813910
  when "110010100110"=> s <="000001000010"; -- Argumento 3238 Funcion -0.96775384
  when "110010100111"=> s <="000001000010"; -- Argumento 3239 Funcion -0.96736629
  when "110010101000"=> s <="000001000011"; -- Argumento 3240 Funcion -0.96697647
  when "110010101001"=> s <="000001000100"; -- Argumento 3241 Funcion -0.96658437
  when "110010101010"=> s <="000001000101"; -- Argumento 3242 Funcion -0.96619000
  when "110010101011"=> s <="000001000110"; -- Argumento 3243 Funcion -0.96579336
  when "110010101100"=> s <="000001000110"; -- Argumento 3244 Funcion -0.96539444
  when "110010101101"=> s <="000001000111"; -- Argumento 3245 Funcion -0.96499325
  when "110010101110"=> s <="000001001000"; -- Argumento 3246 Funcion -0.96458979
  when "110010101111"=> s <="000001001001"; -- Argumento 3247 Funcion -0.96418406
  when "110010110000"=> s <="000001001010"; -- Argumento 3248 Funcion -0.96377607
  when "110010110001"=> s <="000001001011"; -- Argumento 3249 Funcion -0.96336580
  when "110010110010"=> s <="000001001011"; -- Argumento 3250 Funcion -0.96295327
  when "110010110011"=> s <="000001001100"; -- Argumento 3251 Funcion -0.96253847
  when "110010110100"=> s <="000001001101"; -- Argumento 3252 Funcion -0.96212140
  when "110010110101"=> s <="000001001110"; -- Argumento 3253 Funcion -0.96170208
  when "110010110110"=> s <="000001001111"; -- Argumento 3254 Funcion -0.96128049
  when "110010110111"=> s <="000001010000"; -- Argumento 3255 Funcion -0.96085663
  when "110010111000"=> s <="000001010001"; -- Argumento 3256 Funcion -0.96043052
  when "110010111001"=> s <="000001010001"; -- Argumento 3257 Funcion -0.96000215
  when "110010111010"=> s <="000001010010"; -- Argumento 3258 Funcion -0.95957151
  when "110010111011"=> s <="000001010011"; -- Argumento 3259 Funcion -0.95913862
  when "110010111100"=> s <="000001010100"; -- Argumento 3260 Funcion -0.95870347
  when "110010111101"=> s <="000001010101"; -- Argumento 3261 Funcion -0.95826607
  when "110010111110"=> s <="000001010110"; -- Argumento 3262 Funcion -0.95782641
  when "110010111111"=> s <="000001010111"; -- Argumento 3263 Funcion -0.95738450
  when "110011000000"=> s <="000001011000"; -- Argumento 3264 Funcion -0.95694034
  when "110011000001"=> s <="000001011001"; -- Argumento 3265 Funcion -0.95649392
  when "110011000010"=> s <="000001011010"; -- Argumento 3266 Funcion -0.95604525
  when "110011000011"=> s <="000001011010"; -- Argumento 3267 Funcion -0.95559433
  when "110011000100"=> s <="000001011011"; -- Argumento 3268 Funcion -0.95514117
  when "110011000101"=> s <="000001011100"; -- Argumento 3269 Funcion -0.95468575
  when "110011000110"=> s <="000001011101"; -- Argumento 3270 Funcion -0.95422810
  when "110011000111"=> s <="000001011110"; -- Argumento 3271 Funcion -0.95376819
  when "110011001000"=> s <="000001011111"; -- Argumento 3272 Funcion -0.95330604
  when "110011001001"=> s <="000001100000"; -- Argumento 3273 Funcion -0.95284165
  when "110011001010"=> s <="000001100001"; -- Argumento 3274 Funcion -0.95237501
  when "110011001011"=> s <="000001100010"; -- Argumento 3275 Funcion -0.95190614
  when "110011001100"=> s <="000001100011"; -- Argumento 3276 Funcion -0.95143502
  when "110011001101"=> s <="000001100100"; -- Argumento 3277 Funcion -0.95096167
  when "110011001110"=> s <="000001100101"; -- Argumento 3278 Funcion -0.95048607
  when "110011001111"=> s <="000001100110"; -- Argumento 3279 Funcion -0.95000825
  when "110011010000"=> s <="000001100111"; -- Argumento 3280 Funcion -0.94952818
  when "110011010001"=> s <="000001101000"; -- Argumento 3281 Funcion -0.94904588
  when "110011010010"=> s <="000001101001"; -- Argumento 3282 Funcion -0.94856135
  when "110011010011"=> s <="000001101010"; -- Argumento 3283 Funcion -0.94807459
  when "110011010100"=> s <="000001101011"; -- Argumento 3284 Funcion -0.94758559
  when "110011010101"=> s <="000001101100"; -- Argumento 3285 Funcion -0.94709437
  when "110011010110"=> s <="000001101101"; -- Argumento 3286 Funcion -0.94660091
  when "110011010111"=> s <="000001101110"; -- Argumento 3287 Funcion -0.94610523
  when "110011011000"=> s <="000001101111"; -- Argumento 3288 Funcion -0.94560733
  when "110011011001"=> s <="000001110000"; -- Argumento 3289 Funcion -0.94510719
  when "110011011010"=> s <="000001110001"; -- Argumento 3290 Funcion -0.94460484
  when "110011011011"=> s <="000001110010"; -- Argumento 3291 Funcion -0.94410026
  when "110011011100"=> s <="000001110011"; -- Argumento 3292 Funcion -0.94359346
  when "110011011101"=> s <="000001110100"; -- Argumento 3293 Funcion -0.94308444
  when "110011011110"=> s <="000001110101"; -- Argumento 3294 Funcion -0.94257320
  when "110011011111"=> s <="000001110110"; -- Argumento 3295 Funcion -0.94205974
  when "110011100000"=> s <="000001110111"; -- Argumento 3296 Funcion -0.94154407
  when "110011100001"=> s <="000001111000"; -- Argumento 3297 Funcion -0.94102618
  when "110011100010"=> s <="000001111001"; -- Argumento 3298 Funcion -0.94050607
  when "110011100011"=> s <="000001111010"; -- Argumento 3299 Funcion -0.93998375
  when "110011100100"=> s <="000001111011"; -- Argumento 3300 Funcion -0.93945922
  when "110011100101"=> s <="000001111101"; -- Argumento 3301 Funcion -0.93893248
  when "110011100110"=> s <="000001111110"; -- Argumento 3302 Funcion -0.93840353
  when "110011100111"=> s <="000001111111"; -- Argumento 3303 Funcion -0.93787238
  when "110011101000"=> s <="000010000000"; -- Argumento 3304 Funcion -0.93733901
  when "110011101001"=> s <="000010000001"; -- Argumento 3305 Funcion -0.93680344
  when "110011101010"=> s <="000010000010"; -- Argumento 3306 Funcion -0.93626567
  when "110011101011"=> s <="000010000011"; -- Argumento 3307 Funcion -0.93572569
  when "110011101100"=> s <="000010000100"; -- Argumento 3308 Funcion -0.93518351
  when "110011101101"=> s <="000010000101"; -- Argumento 3309 Funcion -0.93463913
  when "110011101110"=> s <="000010000110"; -- Argumento 3310 Funcion -0.93409255
  when "110011101111"=> s <="000010001000"; -- Argumento 3311 Funcion -0.93354377
  when "110011110000"=> s <="000010001001"; -- Argumento 3312 Funcion -0.93299280
  when "110011110001"=> s <="000010001010"; -- Argumento 3313 Funcion -0.93243963
  when "110011110010"=> s <="000010001011"; -- Argumento 3314 Funcion -0.93188427
  when "110011110011"=> s <="000010001100"; -- Argumento 3315 Funcion -0.93132671
  when "110011110100"=> s <="000010001101"; -- Argumento 3316 Funcion -0.93076696
  when "110011110101"=> s <="000010001110"; -- Argumento 3317 Funcion -0.93020502
  when "110011110110"=> s <="000010010000"; -- Argumento 3318 Funcion -0.92964090
  when "110011110111"=> s <="000010010001"; -- Argumento 3319 Funcion -0.92907458
  when "110011111000"=> s <="000010010010"; -- Argumento 3320 Funcion -0.92850608
  when "110011111001"=> s <="000010010011"; -- Argumento 3321 Funcion -0.92793539
  when "110011111010"=> s <="000010010100"; -- Argumento 3322 Funcion -0.92736253
  when "110011111011"=> s <="000010010101"; -- Argumento 3323 Funcion -0.92678747
  when "110011111100"=> s <="000010010111"; -- Argumento 3324 Funcion -0.92621024
  when "110011111101"=> s <="000010011000"; -- Argumento 3325 Funcion -0.92563083
  when "110011111110"=> s <="000010011001"; -- Argumento 3326 Funcion -0.92504924
  when "110011111111"=> s <="000010011010"; -- Argumento 3327 Funcion -0.92446547
  when "110100000000"=> s <="000010011011"; -- Argumento 3328 Funcion -0.92387953
  when "110100000001"=> s <="000010011101"; -- Argumento 3329 Funcion -0.92329142
  when "110100000010"=> s <="000010011110"; -- Argumento 3330 Funcion -0.92270113
  when "110100000011"=> s <="000010011111"; -- Argumento 3331 Funcion -0.92210867
  when "110100000100"=> s <="000010100000"; -- Argumento 3332 Funcion -0.92151404
  when "110100000101"=> s <="000010100001"; -- Argumento 3333 Funcion -0.92091724
  when "110100000110"=> s <="000010100011"; -- Argumento 3334 Funcion -0.92031828
  when "110100000111"=> s <="000010100100"; -- Argumento 3335 Funcion -0.91971715
  when "110100001000"=> s <="000010100101"; -- Argumento 3336 Funcion -0.91911385
  when "110100001001"=> s <="000010100110"; -- Argumento 3337 Funcion -0.91850839
  when "110100001010"=> s <="000010101000"; -- Argumento 3338 Funcion -0.91790078
  when "110100001011"=> s <="000010101001"; -- Argumento 3339 Funcion -0.91729100
  when "110100001100"=> s <="000010101010"; -- Argumento 3340 Funcion -0.91667906
  when "110100001101"=> s <="000010101011"; -- Argumento 3341 Funcion -0.91606497
  when "110100001110"=> s <="000010101101"; -- Argumento 3342 Funcion -0.91544872
  when "110100001111"=> s <="000010101110"; -- Argumento 3343 Funcion -0.91483031
  when "110100010000"=> s <="000010101111"; -- Argumento 3344 Funcion -0.91420976
  when "110100010001"=> s <="000010110000"; -- Argumento 3345 Funcion -0.91358705
  when "110100010010"=> s <="000010110010"; -- Argumento 3346 Funcion -0.91296219
  when "110100010011"=> s <="000010110011"; -- Argumento 3347 Funcion -0.91233518
  when "110100010100"=> s <="000010110100"; -- Argumento 3348 Funcion -0.91170603
  when "110100010101"=> s <="000010110110"; -- Argumento 3349 Funcion -0.91107473
  when "110100010110"=> s <="000010110111"; -- Argumento 3350 Funcion -0.91044129
  when "110100010111"=> s <="000010111000"; -- Argumento 3351 Funcion -0.90980571
  when "110100011000"=> s <="000010111010"; -- Argumento 3352 Funcion -0.90916798
  when "110100011001"=> s <="000010111011"; -- Argumento 3353 Funcion -0.90852812
  when "110100011010"=> s <="000010111100"; -- Argumento 3354 Funcion -0.90788612
  when "110100011011"=> s <="000010111101"; -- Argumento 3355 Funcion -0.90724198
  when "110100011100"=> s <="000010111111"; -- Argumento 3356 Funcion -0.90659570
  when "110100011101"=> s <="000011000000"; -- Argumento 3357 Funcion -0.90594730
  when "110100011110"=> s <="000011000001"; -- Argumento 3358 Funcion -0.90529676
  when "110100011111"=> s <="000011000011"; -- Argumento 3359 Funcion -0.90464409
  when "110100100000"=> s <="000011000100"; -- Argumento 3360 Funcion -0.90398929
  when "110100100001"=> s <="000011000101"; -- Argumento 3361 Funcion -0.90333237
  when "110100100010"=> s <="000011000111"; -- Argumento 3362 Funcion -0.90267332
  when "110100100011"=> s <="000011001000"; -- Argumento 3363 Funcion -0.90201214
  when "110100100100"=> s <="000011001010"; -- Argumento 3364 Funcion -0.90134885
  when "110100100101"=> s <="000011001011"; -- Argumento 3365 Funcion -0.90068343
  when "110100100110"=> s <="000011001100"; -- Argumento 3366 Funcion -0.90001589
  when "110100100111"=> s <="000011001110"; -- Argumento 3367 Funcion -0.89934624
  when "110100101000"=> s <="000011001111"; -- Argumento 3368 Funcion -0.89867447
  when "110100101001"=> s <="000011010000"; -- Argumento 3369 Funcion -0.89800058
  when "110100101010"=> s <="000011010010"; -- Argumento 3370 Funcion -0.89732458
  when "110100101011"=> s <="000011010011"; -- Argumento 3371 Funcion -0.89664647
  when "110100101100"=> s <="000011010101"; -- Argumento 3372 Funcion -0.89596625
  when "110100101101"=> s <="000011010110"; -- Argumento 3373 Funcion -0.89528392
  when "110100101110"=> s <="000011010111"; -- Argumento 3374 Funcion -0.89459949
  when "110100101111"=> s <="000011011001"; -- Argumento 3375 Funcion -0.89391295
  when "110100110000"=> s <="000011011010"; -- Argumento 3376 Funcion -0.89322430
  when "110100110001"=> s <="000011011100"; -- Argumento 3377 Funcion -0.89253356
  when "110100110010"=> s <="000011011101"; -- Argumento 3378 Funcion -0.89184071
  when "110100110011"=> s <="000011011110"; -- Argumento 3379 Funcion -0.89114576
  when "110100110100"=> s <="000011100000"; -- Argumento 3380 Funcion -0.89044872
  when "110100110101"=> s <="000011100001"; -- Argumento 3381 Funcion -0.88974959
  when "110100110110"=> s <="000011100011"; -- Argumento 3382 Funcion -0.88904836
  when "110100110111"=> s <="000011100100"; -- Argumento 3383 Funcion -0.88834503
  when "110100111000"=> s <="000011100110"; -- Argumento 3384 Funcion -0.88763962
  when "110100111001"=> s <="000011100111"; -- Argumento 3385 Funcion -0.88693212
  when "110100111010"=> s <="000011101001"; -- Argumento 3386 Funcion -0.88622253
  when "110100111011"=> s <="000011101010"; -- Argumento 3387 Funcion -0.88551086
  when "110100111100"=> s <="000011101011"; -- Argumento 3388 Funcion -0.88479710
  when "110100111101"=> s <="000011101101"; -- Argumento 3389 Funcion -0.88408126
  when "110100111110"=> s <="000011101110"; -- Argumento 3390 Funcion -0.88336334
  when "110100111111"=> s <="000011110000"; -- Argumento 3391 Funcion -0.88264334
  when "110101000000"=> s <="000011110001"; -- Argumento 3392 Funcion -0.88192126
  when "110101000001"=> s <="000011110011"; -- Argumento 3393 Funcion -0.88119711
  when "110101000010"=> s <="000011110100"; -- Argumento 3394 Funcion -0.88047089
  when "110101000011"=> s <="000011110110"; -- Argumento 3395 Funcion -0.87974259
  when "110101000100"=> s <="000011110111"; -- Argumento 3396 Funcion -0.87901223
  when "110101000101"=> s <="000011111001"; -- Argumento 3397 Funcion -0.87827979
  when "110101000110"=> s <="000011111010"; -- Argumento 3398 Funcion -0.87754529
  when "110101000111"=> s <="000011111100"; -- Argumento 3399 Funcion -0.87680872
  when "110101001000"=> s <="000011111101"; -- Argumento 3400 Funcion -0.87607009
  when "110101001001"=> s <="000011111111"; -- Argumento 3401 Funcion -0.87532940
  when "110101001010"=> s <="000100000000"; -- Argumento 3402 Funcion -0.87458665
  when "110101001011"=> s <="000100000010"; -- Argumento 3403 Funcion -0.87384184
  when "110101001100"=> s <="000100000011"; -- Argumento 3404 Funcion -0.87309498
  when "110101001101"=> s <="000100000101"; -- Argumento 3405 Funcion -0.87234606
  when "110101001110"=> s <="000100000110"; -- Argumento 3406 Funcion -0.87159509
  when "110101001111"=> s <="000100001000"; -- Argumento 3407 Funcion -0.87084206
  when "110101010000"=> s <="000100001010"; -- Argumento 3408 Funcion -0.87008699
  when "110101010001"=> s <="000100001011"; -- Argumento 3409 Funcion -0.86932987
  when "110101010010"=> s <="000100001101"; -- Argumento 3410 Funcion -0.86857071
  when "110101010011"=> s <="000100001110"; -- Argumento 3411 Funcion -0.86780950
  when "110101010100"=> s <="000100010000"; -- Argumento 3412 Funcion -0.86704625
  when "110101010101"=> s <="000100010001"; -- Argumento 3413 Funcion -0.86628095
  when "110101010110"=> s <="000100010011"; -- Argumento 3414 Funcion -0.86551362
  when "110101010111"=> s <="000100010101"; -- Argumento 3415 Funcion -0.86474426
  when "110101011000"=> s <="000100010110"; -- Argumento 3416 Funcion -0.86397286
  when "110101011001"=> s <="000100011000"; -- Argumento 3417 Funcion -0.86319942
  when "110101011010"=> s <="000100011001"; -- Argumento 3418 Funcion -0.86242396
  when "110101011011"=> s <="000100011011"; -- Argumento 3419 Funcion -0.86164646
  when "110101011100"=> s <="000100011100"; -- Argumento 3420 Funcion -0.86086694
  when "110101011101"=> s <="000100011110"; -- Argumento 3421 Funcion -0.86008539
  when "110101011110"=> s <="000100100000"; -- Argumento 3422 Funcion -0.85930182
  when "110101011111"=> s <="000100100001"; -- Argumento 3423 Funcion -0.85851622
  when "110101100000"=> s <="000100100011"; -- Argumento 3424 Funcion -0.85772861
  when "110101100001"=> s <="000100100100"; -- Argumento 3425 Funcion -0.85693898
  when "110101100010"=> s <="000100100110"; -- Argumento 3426 Funcion -0.85614733
  when "110101100011"=> s <="000100101000"; -- Argumento 3427 Funcion -0.85535366
  when "110101100100"=> s <="000100101001"; -- Argumento 3428 Funcion -0.85455799
  when "110101100101"=> s <="000100101011"; -- Argumento 3429 Funcion -0.85376030
  when "110101100110"=> s <="000100101101"; -- Argumento 3430 Funcion -0.85296060
  when "110101100111"=> s <="000100101110"; -- Argumento 3431 Funcion -0.85215890
  when "110101101000"=> s <="000100110000"; -- Argumento 3432 Funcion -0.85135519
  when "110101101001"=> s <="000100110010"; -- Argumento 3433 Funcion -0.85054948
  when "110101101010"=> s <="000100110011"; -- Argumento 3434 Funcion -0.84974177
  when "110101101011"=> s <="000100110101"; -- Argumento 3435 Funcion -0.84893206
  when "110101101100"=> s <="000100110111"; -- Argumento 3436 Funcion -0.84812034
  when "110101101101"=> s <="000100111000"; -- Argumento 3437 Funcion -0.84730664
  when "110101101110"=> s <="000100111010"; -- Argumento 3438 Funcion -0.84649094
  when "110101101111"=> s <="000100111100"; -- Argumento 3439 Funcion -0.84567325
  when "110101110000"=> s <="000100111101"; -- Argumento 3440 Funcion -0.84485357
  when "110101110001"=> s <="000100111111"; -- Argumento 3441 Funcion -0.84403190
  when "110101110010"=> s <="000101000001"; -- Argumento 3442 Funcion -0.84320824
  when "110101110011"=> s <="000101000010"; -- Argumento 3443 Funcion -0.84238260
  when "110101110100"=> s <="000101000100"; -- Argumento 3444 Funcion -0.84155498
  when "110101110101"=> s <="000101000110"; -- Argumento 3445 Funcion -0.84072537
  when "110101110110"=> s <="000101000111"; -- Argumento 3446 Funcion -0.83989379
  when "110101110111"=> s <="000101001001"; -- Argumento 3447 Funcion -0.83906024
  when "110101111000"=> s <="000101001011"; -- Argumento 3448 Funcion -0.83822471
  when "110101111001"=> s <="000101001101"; -- Argumento 3449 Funcion -0.83738720
  when "110101111010"=> s <="000101001110"; -- Argumento 3450 Funcion -0.83654773
  when "110101111011"=> s <="000101010000"; -- Argumento 3451 Funcion -0.83570628
  when "110101111100"=> s <="000101010010"; -- Argumento 3452 Funcion -0.83486287
  when "110101111101"=> s <="000101010011"; -- Argumento 3453 Funcion -0.83401750
  when "110101111110"=> s <="000101010101"; -- Argumento 3454 Funcion -0.83317016
  when "110101111111"=> s <="000101010111"; -- Argumento 3455 Funcion -0.83232087
  when "110110000000"=> s <="000101011001"; -- Argumento 3456 Funcion -0.83146961
  when "110110000001"=> s <="000101011010"; -- Argumento 3457 Funcion -0.83061640
  when "110110000010"=> s <="000101011100"; -- Argumento 3458 Funcion -0.82976123
  when "110110000011"=> s <="000101011110"; -- Argumento 3459 Funcion -0.82890411
  when "110110000100"=> s <="000101100000"; -- Argumento 3460 Funcion -0.82804505
  when "110110000101"=> s <="000101100001"; -- Argumento 3461 Funcion -0.82718403
  when "110110000110"=> s <="000101100011"; -- Argumento 3462 Funcion -0.82632106
  when "110110000111"=> s <="000101100101"; -- Argumento 3463 Funcion -0.82545615
  when "110110001000"=> s <="000101100111"; -- Argumento 3464 Funcion -0.82458930
  when "110110001001"=> s <="000101101001"; -- Argumento 3465 Funcion -0.82372051
  when "110110001010"=> s <="000101101010"; -- Argumento 3466 Funcion -0.82284978
  when "110110001011"=> s <="000101101100"; -- Argumento 3467 Funcion -0.82197712
  when "110110001100"=> s <="000101101110"; -- Argumento 3468 Funcion -0.82110251
  when "110110001101"=> s <="000101110000"; -- Argumento 3469 Funcion -0.82022598
  when "110110001110"=> s <="000101110001"; -- Argumento 3470 Funcion -0.81934752
  when "110110001111"=> s <="000101110011"; -- Argumento 3471 Funcion -0.81846713
  when "110110010000"=> s <="000101110101"; -- Argumento 3472 Funcion -0.81758481
  when "110110010001"=> s <="000101110111"; -- Argumento 3473 Funcion -0.81670057
  when "110110010010"=> s <="000101111001"; -- Argumento 3474 Funcion -0.81581441
  when "110110010011"=> s <="000101111011"; -- Argumento 3475 Funcion -0.81492633
  when "110110010100"=> s <="000101111100"; -- Argumento 3476 Funcion -0.81403633
  when "110110010101"=> s <="000101111110"; -- Argumento 3477 Funcion -0.81314441
  when "110110010110"=> s <="000110000000"; -- Argumento 3478 Funcion -0.81225059
  when "110110010111"=> s <="000110000010"; -- Argumento 3479 Funcion -0.81135485
  when "110110011000"=> s <="000110000100"; -- Argumento 3480 Funcion -0.81045720
  when "110110011001"=> s <="000110000110"; -- Argumento 3481 Funcion -0.80955764
  when "110110011010"=> s <="000110000111"; -- Argumento 3482 Funcion -0.80865618
  when "110110011011"=> s <="000110001001"; -- Argumento 3483 Funcion -0.80775282
  when "110110011100"=> s <="000110001011"; -- Argumento 3484 Funcion -0.80684755
  when "110110011101"=> s <="000110001101"; -- Argumento 3485 Funcion -0.80594039
  when "110110011110"=> s <="000110001111"; -- Argumento 3486 Funcion -0.80503133
  when "110110011111"=> s <="000110010001"; -- Argumento 3487 Funcion -0.80412038
  when "110110100000"=> s <="000110010011"; -- Argumento 3488 Funcion -0.80320753
  when "110110100001"=> s <="000110010100"; -- Argumento 3489 Funcion -0.80229280
  when "110110100010"=> s <="000110010110"; -- Argumento 3490 Funcion -0.80137617
  when "110110100011"=> s <="000110011000"; -- Argumento 3491 Funcion -0.80045766
  when "110110100100"=> s <="000110011010"; -- Argumento 3492 Funcion -0.79953727
  when "110110100101"=> s <="000110011100"; -- Argumento 3493 Funcion -0.79861499
  when "110110100110"=> s <="000110011110"; -- Argumento 3494 Funcion -0.79769084
  when "110110100111"=> s <="000110100000"; -- Argumento 3495 Funcion -0.79676481
  when "110110101000"=> s <="000110100010"; -- Argumento 3496 Funcion -0.79583690
  when "110110101001"=> s <="000110100100"; -- Argumento 3497 Funcion -0.79490713
  when "110110101010"=> s <="000110100101"; -- Argumento 3498 Funcion -0.79397548
  when "110110101011"=> s <="000110100111"; -- Argumento 3499 Funcion -0.79304196
  when "110110101100"=> s <="000110101001"; -- Argumento 3500 Funcion -0.79210658
  when "110110101101"=> s <="000110101011"; -- Argumento 3501 Funcion -0.79116933
  when "110110101110"=> s <="000110101101"; -- Argumento 3502 Funcion -0.79023022
  when "110110101111"=> s <="000110101111"; -- Argumento 3503 Funcion -0.78928925
  when "110110110000"=> s <="000110110001"; -- Argumento 3504 Funcion -0.78834643
  when "110110110001"=> s <="000110110011"; -- Argumento 3505 Funcion -0.78740175
  when "110110110010"=> s <="000110110101"; -- Argumento 3506 Funcion -0.78645521
  when "110110110011"=> s <="000110110111"; -- Argumento 3507 Funcion -0.78550683
  when "110110110100"=> s <="000110111001"; -- Argumento 3508 Funcion -0.78455660
  when "110110110101"=> s <="000110111011"; -- Argumento 3509 Funcion -0.78360452
  when "110110110110"=> s <="000110111101"; -- Argumento 3510 Funcion -0.78265060
  when "110110110111"=> s <="000110111111"; -- Argumento 3511 Funcion -0.78169483
  when "110110111000"=> s <="000111000001"; -- Argumento 3512 Funcion -0.78073723
  when "110110111001"=> s <="000111000011"; -- Argumento 3513 Funcion -0.77977779
  when "110110111010"=> s <="000111000100"; -- Argumento 3514 Funcion -0.77881651
  when "110110111011"=> s <="000111000110"; -- Argumento 3515 Funcion -0.77785340
  when "110110111100"=> s <="000111001000"; -- Argumento 3516 Funcion -0.77688847
  when "110110111101"=> s <="000111001010"; -- Argumento 3517 Funcion -0.77592170
  when "110110111110"=> s <="000111001100"; -- Argumento 3518 Funcion -0.77495311
  when "110110111111"=> s <="000111001110"; -- Argumento 3519 Funcion -0.77398269
  when "110111000000"=> s <="000111010000"; -- Argumento 3520 Funcion -0.77301045
  when "110111000001"=> s <="000111010010"; -- Argumento 3521 Funcion -0.77203640
  when "110111000010"=> s <="000111010100"; -- Argumento 3522 Funcion -0.77106052
  when "110111000011"=> s <="000111010110"; -- Argumento 3523 Funcion -0.77008284
  when "110111000100"=> s <="000111011000"; -- Argumento 3524 Funcion -0.76910334
  when "110111000101"=> s <="000111011010"; -- Argumento 3525 Funcion -0.76812203
  when "110111000110"=> s <="000111011100"; -- Argumento 3526 Funcion -0.76713891
  when "110111000111"=> s <="000111011110"; -- Argumento 3527 Funcion -0.76615399
  when "110111001000"=> s <="000111100000"; -- Argumento 3528 Funcion -0.76516727
  when "110111001001"=> s <="000111100010"; -- Argumento 3529 Funcion -0.76417874
  when "110111001010"=> s <="000111100100"; -- Argumento 3530 Funcion -0.76318842
  when "110111001011"=> s <="000111100111"; -- Argumento 3531 Funcion -0.76219630
  when "110111001100"=> s <="000111101001"; -- Argumento 3532 Funcion -0.76120239
  when "110111001101"=> s <="000111101011"; -- Argumento 3533 Funcion -0.76020668
  when "110111001110"=> s <="000111101101"; -- Argumento 3534 Funcion -0.75920919
  when "110111001111"=> s <="000111101111"; -- Argumento 3535 Funcion -0.75820991
  when "110111010000"=> s <="000111110001"; -- Argumento 3536 Funcion -0.75720885
  when "110111010001"=> s <="000111110011"; -- Argumento 3537 Funcion -0.75620600
  when "110111010010"=> s <="000111110101"; -- Argumento 3538 Funcion -0.75520138
  when "110111010011"=> s <="000111110111"; -- Argumento 3539 Funcion -0.75419498
  when "110111010100"=> s <="000111111001"; -- Argumento 3540 Funcion -0.75318680
  when "110111010101"=> s <="000111111011"; -- Argumento 3541 Funcion -0.75217685
  when "110111010110"=> s <="000111111101"; -- Argumento 3542 Funcion -0.75116513
  when "110111010111"=> s <="000111111111"; -- Argumento 3543 Funcion -0.75015165
  when "110111011000"=> s <="001000000001"; -- Argumento 3544 Funcion -0.74913639
  when "110111011001"=> s <="001000000011"; -- Argumento 3545 Funcion -0.74811938
  when "110111011010"=> s <="001000000101"; -- Argumento 3546 Funcion -0.74710061
  when "110111011011"=> s <="001000001000"; -- Argumento 3547 Funcion -0.74608007
  when "110111011100"=> s <="001000001010"; -- Argumento 3548 Funcion -0.74505779
  when "110111011101"=> s <="001000001100"; -- Argumento 3549 Funcion -0.74403374
  when "110111011110"=> s <="001000001110"; -- Argumento 3550 Funcion -0.74300795
  when "110111011111"=> s <="001000010000"; -- Argumento 3551 Funcion -0.74198041
  when "110111100000"=> s <="001000010010"; -- Argumento 3552 Funcion -0.74095113
  when "110111100001"=> s <="001000010100"; -- Argumento 3553 Funcion -0.73992010
  when "110111100010"=> s <="001000010110"; -- Argumento 3554 Funcion -0.73888732
  when "110111100011"=> s <="001000011000"; -- Argumento 3555 Funcion -0.73785281
  when "110111100100"=> s <="001000011010"; -- Argumento 3556 Funcion -0.73681657
  when "110111100101"=> s <="001000011101"; -- Argumento 3557 Funcion -0.73577859
  when "110111100110"=> s <="001000011111"; -- Argumento 3558 Funcion -0.73473888
  when "110111100111"=> s <="001000100001"; -- Argumento 3559 Funcion -0.73369744
  when "110111101000"=> s <="001000100011"; -- Argumento 3560 Funcion -0.73265427
  when "110111101001"=> s <="001000100101"; -- Argumento 3561 Funcion -0.73160938
  when "110111101010"=> s <="001000100111"; -- Argumento 3562 Funcion -0.73056277
  when "110111101011"=> s <="001000101001"; -- Argumento 3563 Funcion -0.72951444
  when "110111101100"=> s <="001000101100"; -- Argumento 3564 Funcion -0.72846439
  when "110111101101"=> s <="001000101110"; -- Argumento 3565 Funcion -0.72741263
  when "110111101110"=> s <="001000110000"; -- Argumento 3566 Funcion -0.72635916
  when "110111101111"=> s <="001000110010"; -- Argumento 3567 Funcion -0.72530397
  when "110111110000"=> s <="001000110100"; -- Argumento 3568 Funcion -0.72424708
  when "110111110001"=> s <="001000110110"; -- Argumento 3569 Funcion -0.72318849
  when "110111110010"=> s <="001000111001"; -- Argumento 3570 Funcion -0.72212819
  when "110111110011"=> s <="001000111011"; -- Argumento 3571 Funcion -0.72106620
  when "110111110100"=> s <="001000111101"; -- Argumento 3572 Funcion -0.72000251
  when "110111110101"=> s <="001000111111"; -- Argumento 3573 Funcion -0.71893712
  when "110111110110"=> s <="001001000001"; -- Argumento 3574 Funcion -0.71787005
  when "110111110111"=> s <="001001000011"; -- Argumento 3575 Funcion -0.71680128
  when "110111111000"=> s <="001001000110"; -- Argumento 3576 Funcion -0.71573083
  when "110111111001"=> s <="001001001000"; -- Argumento 3577 Funcion -0.71465869
  when "110111111010"=> s <="001001001010"; -- Argumento 3578 Funcion -0.71358487
  when "110111111011"=> s <="001001001100"; -- Argumento 3579 Funcion -0.71250937
  when "110111111100"=> s <="001001001110"; -- Argumento 3580 Funcion -0.71143220
  when "110111111101"=> s <="001001010001"; -- Argumento 3581 Funcion -0.71035335
  when "110111111110"=> s <="001001010011"; -- Argumento 3582 Funcion -0.70927283
  when "110111111111"=> s <="001001010101"; -- Argumento 3583 Funcion -0.70819064
  when "111000000000"=> s <="001001010111"; -- Argumento 3584 Funcion -0.70710678
  when "111000000001"=> s <="001001011010"; -- Argumento 3585 Funcion -0.70602126
  when "111000000010"=> s <="001001011100"; -- Argumento 3586 Funcion -0.70493408
  when "111000000011"=> s <="001001011110"; -- Argumento 3587 Funcion -0.70384524
  when "111000000100"=> s <="001001100000"; -- Argumento 3588 Funcion -0.70275474
  when "111000000101"=> s <="001001100010"; -- Argumento 3589 Funcion -0.70166259
  when "111000000110"=> s <="001001100101"; -- Argumento 3590 Funcion -0.70056879
  when "111000000111"=> s <="001001100111"; -- Argumento 3591 Funcion -0.69947334
  when "111000001000"=> s <="001001101001"; -- Argumento 3592 Funcion -0.69837625
  when "111000001001"=> s <="001001101011"; -- Argumento 3593 Funcion -0.69727751
  when "111000001010"=> s <="001001101110"; -- Argumento 3594 Funcion -0.69617713
  when "111000001011"=> s <="001001110000"; -- Argumento 3595 Funcion -0.69507511
  when "111000001100"=> s <="001001110010"; -- Argumento 3596 Funcion -0.69397146
  when "111000001101"=> s <="001001110101"; -- Argumento 3597 Funcion -0.69286617
  when "111000001110"=> s <="001001110111"; -- Argumento 3598 Funcion -0.69175926
  when "111000001111"=> s <="001001111001"; -- Argumento 3599 Funcion -0.69065071
  when "111000010000"=> s <="001001111011"; -- Argumento 3600 Funcion -0.68954054
  when "111000010001"=> s <="001001111110"; -- Argumento 3601 Funcion -0.68842875
  when "111000010010"=> s <="001010000000"; -- Argumento 3602 Funcion -0.68731534
  when "111000010011"=> s <="001010000010"; -- Argumento 3603 Funcion -0.68620031
  when "111000010100"=> s <="001010000100"; -- Argumento 3604 Funcion -0.68508367
  when "111000010101"=> s <="001010000111"; -- Argumento 3605 Funcion -0.68396541
  when "111000010110"=> s <="001010001001"; -- Argumento 3606 Funcion -0.68284555
  when "111000010111"=> s <="001010001011"; -- Argumento 3607 Funcion -0.68172407
  when "111000011000"=> s <="001010001110"; -- Argumento 3608 Funcion -0.68060100
  when "111000011001"=> s <="001010010000"; -- Argumento 3609 Funcion -0.67947632
  when "111000011010"=> s <="001010010010"; -- Argumento 3610 Funcion -0.67835004
  when "111000011011"=> s <="001010010101"; -- Argumento 3611 Funcion -0.67722217
  when "111000011100"=> s <="001010010111"; -- Argumento 3612 Funcion -0.67609270
  when "111000011101"=> s <="001010011001"; -- Argumento 3613 Funcion -0.67496165
  when "111000011110"=> s <="001010011011"; -- Argumento 3614 Funcion -0.67382900
  when "111000011111"=> s <="001010011110"; -- Argumento 3615 Funcion -0.67269477
  when "111000100000"=> s <="001010100000"; -- Argumento 3616 Funcion -0.67155895
  when "111000100001"=> s <="001010100010"; -- Argumento 3617 Funcion -0.67042156
  when "111000100010"=> s <="001010100101"; -- Argumento 3618 Funcion -0.66928259
  when "111000100011"=> s <="001010100111"; -- Argumento 3619 Funcion -0.66814204
  when "111000100100"=> s <="001010101001"; -- Argumento 3620 Funcion -0.66699992
  when "111000100101"=> s <="001010101100"; -- Argumento 3621 Funcion -0.66585623
  when "111000100110"=> s <="001010101110"; -- Argumento 3622 Funcion -0.66471098
  when "111000100111"=> s <="001010110001"; -- Argumento 3623 Funcion -0.66356416
  when "111000101000"=> s <="001010110011"; -- Argumento 3624 Funcion -0.66241578
  when "111000101001"=> s <="001010110101"; -- Argumento 3625 Funcion -0.66126584
  when "111000101010"=> s <="001010111000"; -- Argumento 3626 Funcion -0.66011434
  when "111000101011"=> s <="001010111010"; -- Argumento 3627 Funcion -0.65896129
  when "111000101100"=> s <="001010111100"; -- Argumento 3628 Funcion -0.65780669
  when "111000101101"=> s <="001010111111"; -- Argumento 3629 Funcion -0.65665055
  when "111000101110"=> s <="001011000001"; -- Argumento 3630 Funcion -0.65549285
  when "111000101111"=> s <="001011000011"; -- Argumento 3631 Funcion -0.65433362
  when "111000110000"=> s <="001011000110"; -- Argumento 3632 Funcion -0.65317284
  when "111000110001"=> s <="001011001000"; -- Argumento 3633 Funcion -0.65201053
  when "111000110010"=> s <="001011001011"; -- Argumento 3634 Funcion -0.65084668
  when "111000110011"=> s <="001011001101"; -- Argumento 3635 Funcion -0.64968131
  when "111000110100"=> s <="001011001111"; -- Argumento 3636 Funcion -0.64851440
  when "111000110101"=> s <="001011010010"; -- Argumento 3637 Funcion -0.64734597
  when "111000110110"=> s <="001011010100"; -- Argumento 3638 Funcion -0.64617601
  when "111000110111"=> s <="001011010111"; -- Argumento 3639 Funcion -0.64500454
  when "111000111000"=> s <="001011011001"; -- Argumento 3640 Funcion -0.64383154
  when "111000111001"=> s <="001011011011"; -- Argumento 3641 Funcion -0.64265703
  when "111000111010"=> s <="001011011110"; -- Argumento 3642 Funcion -0.64148101
  when "111000111011"=> s <="001011100000"; -- Argumento 3643 Funcion -0.64030348
  when "111000111100"=> s <="001011100011"; -- Argumento 3644 Funcion -0.63912444
  when "111000111101"=> s <="001011100101"; -- Argumento 3645 Funcion -0.63794390
  when "111000111110"=> s <="001011100111"; -- Argumento 3646 Funcion -0.63676186
  when "111000111111"=> s <="001011101010"; -- Argumento 3647 Funcion -0.63557832
  when "111001000000"=> s <="001011101100"; -- Argumento 3648 Funcion -0.63439328
  when "111001000001"=> s <="001011101111"; -- Argumento 3649 Funcion -0.63320676
  when "111001000010"=> s <="001011110001"; -- Argumento 3650 Funcion -0.63201874
  when "111001000011"=> s <="001011110100"; -- Argumento 3651 Funcion -0.63082923
  when "111001000100"=> s <="001011110110"; -- Argumento 3652 Funcion -0.62963824
  when "111001000101"=> s <="001011111000"; -- Argumento 3653 Funcion -0.62844577
  when "111001000110"=> s <="001011111011"; -- Argumento 3654 Funcion -0.62725182
  when "111001000111"=> s <="001011111101"; -- Argumento 3655 Funcion -0.62605639
  when "111001001000"=> s <="001100000000"; -- Argumento 3656 Funcion -0.62485949
  when "111001001001"=> s <="001100000010"; -- Argumento 3657 Funcion -0.62366112
  when "111001001010"=> s <="001100000101"; -- Argumento 3658 Funcion -0.62246128
  when "111001001011"=> s <="001100000111"; -- Argumento 3659 Funcion -0.62125998
  when "111001001100"=> s <="001100001010"; -- Argumento 3660 Funcion -0.62005721
  when "111001001101"=> s <="001100001100"; -- Argumento 3661 Funcion -0.61885299
  when "111001001110"=> s <="001100001111"; -- Argumento 3662 Funcion -0.61764731
  when "111001001111"=> s <="001100010001"; -- Argumento 3663 Funcion -0.61644017
  when "111001010000"=> s <="001100010100"; -- Argumento 3664 Funcion -0.61523159
  when "111001010001"=> s <="001100010110"; -- Argumento 3665 Funcion -0.61402156
  when "111001010010"=> s <="001100011000"; -- Argumento 3666 Funcion -0.61281008
  when "111001010011"=> s <="001100011011"; -- Argumento 3667 Funcion -0.61159716
  when "111001010100"=> s <="001100011101"; -- Argumento 3668 Funcion -0.61038281
  when "111001010101"=> s <="001100100000"; -- Argumento 3669 Funcion -0.60916701
  when "111001010110"=> s <="001100100010"; -- Argumento 3670 Funcion -0.60794978
  when "111001010111"=> s <="001100100101"; -- Argumento 3671 Funcion -0.60673113
  when "111001011000"=> s <="001100100111"; -- Argumento 3672 Funcion -0.60551104
  when "111001011001"=> s <="001100101010"; -- Argumento 3673 Funcion -0.60428953
  when "111001011010"=> s <="001100101100"; -- Argumento 3674 Funcion -0.60306660
  when "111001011011"=> s <="001100101111"; -- Argumento 3675 Funcion -0.60184225
  when "111001011100"=> s <="001100110001"; -- Argumento 3676 Funcion -0.60061648
  when "111001011101"=> s <="001100110100"; -- Argumento 3677 Funcion -0.59938930
  when "111001011110"=> s <="001100110110"; -- Argumento 3678 Funcion -0.59816071
  when "111001011111"=> s <="001100111001"; -- Argumento 3679 Funcion -0.59693071
  when "111001100000"=> s <="001100111100"; -- Argumento 3680 Funcion -0.59569930
  when "111001100001"=> s <="001100111110"; -- Argumento 3681 Funcion -0.59446650
  when "111001100010"=> s <="001101000001"; -- Argumento 3682 Funcion -0.59323230
  when "111001100011"=> s <="001101000011"; -- Argumento 3683 Funcion -0.59199669
  when "111001100100"=> s <="001101000110"; -- Argumento 3684 Funcion -0.59075970
  when "111001100101"=> s <="001101001000"; -- Argumento 3685 Funcion -0.58952132
  when "111001100110"=> s <="001101001011"; -- Argumento 3686 Funcion -0.58828155
  when "111001100111"=> s <="001101001101"; -- Argumento 3687 Funcion -0.58704039
  when "111001101000"=> s <="001101010000"; -- Argumento 3688 Funcion -0.58579786
  when "111001101001"=> s <="001101010010"; -- Argumento 3689 Funcion -0.58455394
  when "111001101010"=> s <="001101010101"; -- Argumento 3690 Funcion -0.58330865
  when "111001101011"=> s <="001101010111"; -- Argumento 3691 Funcion -0.58206199
  when "111001101100"=> s <="001101011010"; -- Argumento 3692 Funcion -0.58081396
  when "111001101101"=> s <="001101011101"; -- Argumento 3693 Funcion -0.57956456
  when "111001101110"=> s <="001101011111"; -- Argumento 3694 Funcion -0.57831380
  when "111001101111"=> s <="001101100010"; -- Argumento 3695 Funcion -0.57706167
  when "111001110000"=> s <="001101100100"; -- Argumento 3696 Funcion -0.57580819
  when "111001110001"=> s <="001101100111"; -- Argumento 3697 Funcion -0.57455336
  when "111001110010"=> s <="001101101001"; -- Argumento 3698 Funcion -0.57329717
  when "111001110011"=> s <="001101101100"; -- Argumento 3699 Funcion -0.57203963
  when "111001110100"=> s <="001101101111"; -- Argumento 3700 Funcion -0.57078075
  when "111001110101"=> s <="001101110001"; -- Argumento 3701 Funcion -0.56952052
  when "111001110110"=> s <="001101110100"; -- Argumento 3702 Funcion -0.56825895
  when "111001110111"=> s <="001101110110"; -- Argumento 3703 Funcion -0.56699605
  when "111001111000"=> s <="001101111001"; -- Argumento 3704 Funcion -0.56573181
  when "111001111001"=> s <="001101111011"; -- Argumento 3705 Funcion -0.56446624
  when "111001111010"=> s <="001101111110"; -- Argumento 3706 Funcion -0.56319934
  when "111001111011"=> s <="001110000001"; -- Argumento 3707 Funcion -0.56193112
  when "111001111100"=> s <="001110000011"; -- Argumento 3708 Funcion -0.56066158
  when "111001111101"=> s <="001110000110"; -- Argumento 3709 Funcion -0.55939071
  when "111001111110"=> s <="001110001000"; -- Argumento 3710 Funcion -0.55811853
  when "111001111111"=> s <="001110001011"; -- Argumento 3711 Funcion -0.55684504
  when "111010000000"=> s <="001110001110"; -- Argumento 3712 Funcion -0.55557023
  when "111010000001"=> s <="001110010000"; -- Argumento 3713 Funcion -0.55429412
  when "111010000010"=> s <="001110010011"; -- Argumento 3714 Funcion -0.55301671
  when "111010000011"=> s <="001110010110"; -- Argumento 3715 Funcion -0.55173799
  when "111010000100"=> s <="001110011000"; -- Argumento 3716 Funcion -0.55045797
  when "111010000101"=> s <="001110011011"; -- Argumento 3717 Funcion -0.54917666
  when "111010000110"=> s <="001110011101"; -- Argumento 3718 Funcion -0.54789406
  when "111010000111"=> s <="001110100000"; -- Argumento 3719 Funcion -0.54661017
  when "111010001000"=> s <="001110100011"; -- Argumento 3720 Funcion -0.54532499
  when "111010001001"=> s <="001110100101"; -- Argumento 3721 Funcion -0.54403853
  when "111010001010"=> s <="001110101000"; -- Argumento 3722 Funcion -0.54275078
  when "111010001011"=> s <="001110101011"; -- Argumento 3723 Funcion -0.54146177
  when "111010001100"=> s <="001110101101"; -- Argumento 3724 Funcion -0.54017147
  when "111010001101"=> s <="001110110000"; -- Argumento 3725 Funcion -0.53887991
  when "111010001110"=> s <="001110110011"; -- Argumento 3726 Funcion -0.53758708
  when "111010001111"=> s <="001110110101"; -- Argumento 3727 Funcion -0.53629298
  when "111010010000"=> s <="001110111000"; -- Argumento 3728 Funcion -0.53499762
  when "111010010001"=> s <="001110111010"; -- Argumento 3729 Funcion -0.53370100
  when "111010010010"=> s <="001110111101"; -- Argumento 3730 Funcion -0.53240313
  when "111010010011"=> s <="001111000000"; -- Argumento 3731 Funcion -0.53110400
  when "111010010100"=> s <="001111000010"; -- Argumento 3732 Funcion -0.52980362
  when "111010010101"=> s <="001111000101"; -- Argumento 3733 Funcion -0.52850200
  when "111010010110"=> s <="001111001000"; -- Argumento 3734 Funcion -0.52719913
  when "111010010111"=> s <="001111001010"; -- Argumento 3735 Funcion -0.52589503
  when "111010011000"=> s <="001111001101"; -- Argumento 3736 Funcion -0.52458968
  when "111010011001"=> s <="001111010000"; -- Argumento 3737 Funcion -0.52328310
  when "111010011010"=> s <="001111010010"; -- Argumento 3738 Funcion -0.52197529
  when "111010011011"=> s <="001111010101"; -- Argumento 3739 Funcion -0.52066625
  when "111010011100"=> s <="001111011000"; -- Argumento 3740 Funcion -0.51935599
  when "111010011101"=> s <="001111011011"; -- Argumento 3741 Funcion -0.51804450
  when "111010011110"=> s <="001111011101"; -- Argumento 3742 Funcion -0.51673180
  when "111010011111"=> s <="001111100000"; -- Argumento 3743 Funcion -0.51541788
  when "111010100000"=> s <="001111100011"; -- Argumento 3744 Funcion -0.51410274
  when "111010100001"=> s <="001111100101"; -- Argumento 3745 Funcion -0.51278640
  when "111010100010"=> s <="001111101000"; -- Argumento 3746 Funcion -0.51146885
  when "111010100011"=> s <="001111101011"; -- Argumento 3747 Funcion -0.51015010
  when "111010100100"=> s <="001111101101"; -- Argumento 3748 Funcion -0.50883014
  when "111010100101"=> s <="001111110000"; -- Argumento 3749 Funcion -0.50750899
  when "111010100110"=> s <="001111110011"; -- Argumento 3750 Funcion -0.50618665
  when "111010100111"=> s <="001111110110"; -- Argumento 3751 Funcion -0.50486311
  when "111010101000"=> s <="001111111000"; -- Argumento 3752 Funcion -0.50353838
  when "111010101001"=> s <="001111111011"; -- Argumento 3753 Funcion -0.50221247
  when "111010101010"=> s <="001111111110"; -- Argumento 3754 Funcion -0.50088538
  when "111010101011"=> s <="010000000000"; -- Argumento 3755 Funcion -0.49955711
  when "111010101100"=> s <="010000000011"; -- Argumento 3756 Funcion -0.49822767
  when "111010101101"=> s <="010000000110"; -- Argumento 3757 Funcion -0.49689705
  when "111010101110"=> s <="010000001001"; -- Argumento 3758 Funcion -0.49556526
  when "111010101111"=> s <="010000001011"; -- Argumento 3759 Funcion -0.49423231
  when "111010110000"=> s <="010000001110"; -- Argumento 3760 Funcion -0.49289819
  when "111010110001"=> s <="010000010001"; -- Argumento 3761 Funcion -0.49156292
  when "111010110010"=> s <="010000010100"; -- Argumento 3762 Funcion -0.49022648
  when "111010110011"=> s <="010000010110"; -- Argumento 3763 Funcion -0.48888890
  when "111010110100"=> s <="010000011001"; -- Argumento 3764 Funcion -0.48755016
  when "111010110101"=> s <="010000011100"; -- Argumento 3765 Funcion -0.48621028
  when "111010110110"=> s <="010000011110"; -- Argumento 3766 Funcion -0.48486925
  when "111010110111"=> s <="010000100001"; -- Argumento 3767 Funcion -0.48352708
  when "111010111000"=> s <="010000100100"; -- Argumento 3768 Funcion -0.48218377
  when "111010111001"=> s <="010000100111"; -- Argumento 3769 Funcion -0.48083933
  when "111010111010"=> s <="010000101001"; -- Argumento 3770 Funcion -0.47949376
  when "111010111011"=> s <="010000101100"; -- Argumento 3771 Funcion -0.47814706
  when "111010111100"=> s <="010000101111"; -- Argumento 3772 Funcion -0.47679923
  when "111010111101"=> s <="010000110010"; -- Argumento 3773 Funcion -0.47545028
  when "111010111110"=> s <="010000110101"; -- Argumento 3774 Funcion -0.47410021
  when "111010111111"=> s <="010000110111"; -- Argumento 3775 Funcion -0.47274903
  when "111011000000"=> s <="010000111010"; -- Argumento 3776 Funcion -0.47139674
  when "111011000001"=> s <="010000111101"; -- Argumento 3777 Funcion -0.47004333
  when "111011000010"=> s <="010001000000"; -- Argumento 3778 Funcion -0.46868882
  when "111011000011"=> s <="010001000010"; -- Argumento 3779 Funcion -0.46733321
  when "111011000100"=> s <="010001000101"; -- Argumento 3780 Funcion -0.46597650
  when "111011000101"=> s <="010001001000"; -- Argumento 3781 Funcion -0.46461869
  when "111011000110"=> s <="010001001011"; -- Argumento 3782 Funcion -0.46325978
  when "111011000111"=> s <="010001001110"; -- Argumento 3783 Funcion -0.46189979
  when "111011001000"=> s <="010001010000"; -- Argumento 3784 Funcion -0.46053871
  when "111011001001"=> s <="010001010011"; -- Argumento 3785 Funcion -0.45917655
  when "111011001010"=> s <="010001010110"; -- Argumento 3786 Funcion -0.45781330
  when "111011001011"=> s <="010001011001"; -- Argumento 3787 Funcion -0.45644898
  when "111011001100"=> s <="010001011011"; -- Argumento 3788 Funcion -0.45508359
  when "111011001101"=> s <="010001011110"; -- Argumento 3789 Funcion -0.45371712
  when "111011001110"=> s <="010001100001"; -- Argumento 3790 Funcion -0.45234959
  when "111011001111"=> s <="010001100100"; -- Argumento 3791 Funcion -0.45098099
  when "111011010000"=> s <="010001100111"; -- Argumento 3792 Funcion -0.44961133
  when "111011010001"=> s <="010001101010"; -- Argumento 3793 Funcion -0.44824061
  when "111011010010"=> s <="010001101100"; -- Argumento 3794 Funcion -0.44686884
  when "111011010011"=> s <="010001101111"; -- Argumento 3795 Funcion -0.44549602
  when "111011010100"=> s <="010001110010"; -- Argumento 3796 Funcion -0.44412214
  when "111011010101"=> s <="010001110101"; -- Argumento 3797 Funcion -0.44274723
  when "111011010110"=> s <="010001111000"; -- Argumento 3798 Funcion -0.44137127
  when "111011010111"=> s <="010001111010"; -- Argumento 3799 Funcion -0.43999427
  when "111011011000"=> s <="010001111101"; -- Argumento 3800 Funcion -0.43861624
  when "111011011001"=> s <="010010000000"; -- Argumento 3801 Funcion -0.43723717
  when "111011011010"=> s <="010010000011"; -- Argumento 3802 Funcion -0.43585708
  when "111011011011"=> s <="010010000110"; -- Argumento 3803 Funcion -0.43447596
  when "111011011100"=> s <="010010001001"; -- Argumento 3804 Funcion -0.43309382
  when "111011011101"=> s <="010010001011"; -- Argumento 3805 Funcion -0.43171066
  when "111011011110"=> s <="010010001110"; -- Argumento 3806 Funcion -0.43032648
  when "111011011111"=> s <="010010010001"; -- Argumento 3807 Funcion -0.42894129
  when "111011100000"=> s <="010010010100"; -- Argumento 3808 Funcion -0.42755509
  when "111011100001"=> s <="010010010111"; -- Argumento 3809 Funcion -0.42616789
  when "111011100010"=> s <="010010011010"; -- Argumento 3810 Funcion -0.42477968
  when "111011100011"=> s <="010010011100"; -- Argumento 3811 Funcion -0.42339047
  when "111011100100"=> s <="010010011111"; -- Argumento 3812 Funcion -0.42200027
  when "111011100101"=> s <="010010100010"; -- Argumento 3813 Funcion -0.42060907
  when "111011100110"=> s <="010010100101"; -- Argumento 3814 Funcion -0.41921689
  when "111011100111"=> s <="010010101000"; -- Argumento 3815 Funcion -0.41782372
  when "111011101000"=> s <="010010101011"; -- Argumento 3816 Funcion -0.41642956
  when "111011101001"=> s <="010010101110"; -- Argumento 3817 Funcion -0.41503442
  when "111011101010"=> s <="010010110000"; -- Argumento 3818 Funcion -0.41363831
  when "111011101011"=> s <="010010110011"; -- Argumento 3819 Funcion -0.41224123
  when "111011101100"=> s <="010010110110"; -- Argumento 3820 Funcion -0.41084317
  when "111011101101"=> s <="010010111001"; -- Argumento 3821 Funcion -0.40944415
  when "111011101110"=> s <="010010111100"; -- Argumento 3822 Funcion -0.40804416
  when "111011101111"=> s <="010010111111"; -- Argumento 3823 Funcion -0.40664322
  when "111011110000"=> s <="010011000010"; -- Argumento 3824 Funcion -0.40524131
  when "111011110001"=> s <="010011000100"; -- Argumento 3825 Funcion -0.40383846
  when "111011110010"=> s <="010011000111"; -- Argumento 3826 Funcion -0.40243465
  when "111011110011"=> s <="010011001010"; -- Argumento 3827 Funcion -0.40102990
  when "111011110100"=> s <="010011001101"; -- Argumento 3828 Funcion -0.39962420
  when "111011110101"=> s <="010011010000"; -- Argumento 3829 Funcion -0.39821756
  when "111011110110"=> s <="010011010011"; -- Argumento 3830 Funcion -0.39680999
  when "111011110111"=> s <="010011010110"; -- Argumento 3831 Funcion -0.39540148
  when "111011111000"=> s <="010011011001"; -- Argumento 3832 Funcion -0.39399204
  when "111011111001"=> s <="010011011011"; -- Argumento 3833 Funcion -0.39258167
  when "111011111010"=> s <="010011011110"; -- Argumento 3834 Funcion -0.39117038
  when "111011111011"=> s <="010011100001"; -- Argumento 3835 Funcion -0.38975817
  when "111011111100"=> s <="010011100100"; -- Argumento 3836 Funcion -0.38834505
  when "111011111101"=> s <="010011100111"; -- Argumento 3837 Funcion -0.38693101
  when "111011111110"=> s <="010011101010"; -- Argumento 3838 Funcion -0.38551605
  when "111011111111"=> s <="010011101101"; -- Argumento 3839 Funcion -0.38410020
  when "111100000000"=> s <="010011110000"; -- Argumento 3840 Funcion -0.38268343
  when "111100000001"=> s <="010011110011"; -- Argumento 3841 Funcion -0.38126577
  when "111100000010"=> s <="010011110110"; -- Argumento 3842 Funcion -0.37984721
  when "111100000011"=> s <="010011111000"; -- Argumento 3843 Funcion -0.37842775
  when "111100000100"=> s <="010011111011"; -- Argumento 3844 Funcion -0.37700741
  when "111100000101"=> s <="010011111110"; -- Argumento 3845 Funcion -0.37558618
  when "111100000110"=> s <="010100000001"; -- Argumento 3846 Funcion -0.37416406
  when "111100000111"=> s <="010100000100"; -- Argumento 3847 Funcion -0.37274107
  when "111100001000"=> s <="010100000111"; -- Argumento 3848 Funcion -0.37131719
  when "111100001001"=> s <="010100001010"; -- Argumento 3849 Funcion -0.36989245
  when "111100001010"=> s <="010100001101"; -- Argumento 3850 Funcion -0.36846683
  when "111100001011"=> s <="010100010000"; -- Argumento 3851 Funcion -0.36704035
  when "111100001100"=> s <="010100010011"; -- Argumento 3852 Funcion -0.36561300
  when "111100001101"=> s <="010100010110"; -- Argumento 3853 Funcion -0.36418479
  when "111100001110"=> s <="010100011001"; -- Argumento 3854 Funcion -0.36275572
  when "111100001111"=> s <="010100011100"; -- Argumento 3855 Funcion -0.36132581
  when "111100010000"=> s <="010100011110"; -- Argumento 3856 Funcion -0.35989504
  when "111100010001"=> s <="010100100001"; -- Argumento 3857 Funcion -0.35846342
  when "111100010010"=> s <="010100100100"; -- Argumento 3858 Funcion -0.35703096
  when "111100010011"=> s <="010100100111"; -- Argumento 3859 Funcion -0.35559766
  when "111100010100"=> s <="010100101010"; -- Argumento 3860 Funcion -0.35416353
  when "111100010101"=> s <="010100101101"; -- Argumento 3861 Funcion -0.35272856
  when "111100010110"=> s <="010100110000"; -- Argumento 3862 Funcion -0.35129276
  when "111100010111"=> s <="010100110011"; -- Argumento 3863 Funcion -0.34985613
  when "111100011000"=> s <="010100110110"; -- Argumento 3864 Funcion -0.34841868
  when "111100011001"=> s <="010100111001"; -- Argumento 3865 Funcion -0.34698041
  when "111100011010"=> s <="010100111100"; -- Argumento 3866 Funcion -0.34554132
  when "111100011011"=> s <="010100111111"; -- Argumento 3867 Funcion -0.34410143
  when "111100011100"=> s <="010101000010"; -- Argumento 3868 Funcion -0.34266072
  when "111100011101"=> s <="010101000101"; -- Argumento 3869 Funcion -0.34121920
  when "111100011110"=> s <="010101001000"; -- Argumento 3870 Funcion -0.33977688
  when "111100011111"=> s <="010101001011"; -- Argumento 3871 Funcion -0.33833377
  when "111100100000"=> s <="010101001110"; -- Argumento 3872 Funcion -0.33688985
  when "111100100001"=> s <="010101010001"; -- Argumento 3873 Funcion -0.33544515
  when "111100100010"=> s <="010101010011"; -- Argumento 3874 Funcion -0.33399965
  when "111100100011"=> s <="010101010110"; -- Argumento 3875 Funcion -0.33255337
  when "111100100100"=> s <="010101011001"; -- Argumento 3876 Funcion -0.33110631
  when "111100100101"=> s <="010101011100"; -- Argumento 3877 Funcion -0.32965846
  when "111100100110"=> s <="010101011111"; -- Argumento 3878 Funcion -0.32820984
  when "111100100111"=> s <="010101100010"; -- Argumento 3879 Funcion -0.32676045
  when "111100101000"=> s <="010101100101"; -- Argumento 3880 Funcion -0.32531029
  when "111100101001"=> s <="010101101000"; -- Argumento 3881 Funcion -0.32385937
  when "111100101010"=> s <="010101101011"; -- Argumento 3882 Funcion -0.32240768
  when "111100101011"=> s <="010101101110"; -- Argumento 3883 Funcion -0.32095523
  when "111100101100"=> s <="010101110001"; -- Argumento 3884 Funcion -0.31950203
  when "111100101101"=> s <="010101110100"; -- Argumento 3885 Funcion -0.31804808
  when "111100101110"=> s <="010101110111"; -- Argumento 3886 Funcion -0.31659338
  when "111100101111"=> s <="010101111010"; -- Argumento 3887 Funcion -0.31513793
  when "111100110000"=> s <="010101111101"; -- Argumento 3888 Funcion -0.31368174
  when "111100110001"=> s <="010110000000"; -- Argumento 3889 Funcion -0.31222481
  when "111100110010"=> s <="010110000011"; -- Argumento 3890 Funcion -0.31076715
  when "111100110011"=> s <="010110000110"; -- Argumento 3891 Funcion -0.30930876
  when "111100110100"=> s <="010110001001"; -- Argumento 3892 Funcion -0.30784964
  when "111100110101"=> s <="010110001100"; -- Argumento 3893 Funcion -0.30638980
  when "111100110110"=> s <="010110001111"; -- Argumento 3894 Funcion -0.30492923
  when "111100110111"=> s <="010110010010"; -- Argumento 3895 Funcion -0.30346795
  when "111100111000"=> s <="010110010101"; -- Argumento 3896 Funcion -0.30200595
  when "111100111001"=> s <="010110011000"; -- Argumento 3897 Funcion -0.30054324
  when "111100111010"=> s <="010110011011"; -- Argumento 3898 Funcion -0.29907983
  when "111100111011"=> s <="010110011110"; -- Argumento 3899 Funcion -0.29761571
  when "111100111100"=> s <="010110100001"; -- Argumento 3900 Funcion -0.29615089
  when "111100111101"=> s <="010110100100"; -- Argumento 3901 Funcion -0.29468537
  when "111100111110"=> s <="010110100111"; -- Argumento 3902 Funcion -0.29321916
  when "111100111111"=> s <="010110101010"; -- Argumento 3903 Funcion -0.29175226
  when "111101000000"=> s <="010110101101"; -- Argumento 3904 Funcion -0.29028468
  when "111101000001"=> s <="010110110000"; -- Argumento 3905 Funcion -0.28881641
  when "111101000010"=> s <="010110110011"; -- Argumento 3906 Funcion -0.28734746
  when "111101000011"=> s <="010110110110"; -- Argumento 3907 Funcion -0.28587783
  when "111101000100"=> s <="010110111001"; -- Argumento 3908 Funcion -0.28440754
  when "111101000101"=> s <="010110111100"; -- Argumento 3909 Funcion -0.28293657
  when "111101000110"=> s <="010110111111"; -- Argumento 3910 Funcion -0.28146494
  when "111101000111"=> s <="010111000010"; -- Argumento 3911 Funcion -0.27999264
  when "111101001000"=> s <="010111000101"; -- Argumento 3912 Funcion -0.27851969
  when "111101001001"=> s <="010111001000"; -- Argumento 3913 Funcion -0.27704608
  when "111101001010"=> s <="010111001011"; -- Argumento 3914 Funcion -0.27557182
  when "111101001011"=> s <="010111001110"; -- Argumento 3915 Funcion -0.27409691
  when "111101001100"=> s <="010111010001"; -- Argumento 3916 Funcion -0.27262136
  when "111101001101"=> s <="010111010100"; -- Argumento 3917 Funcion -0.27114516
  when "111101001110"=> s <="010111010111"; -- Argumento 3918 Funcion -0.26966833
  when "111101001111"=> s <="010111011010"; -- Argumento 3919 Funcion -0.26819086
  when "111101010000"=> s <="010111011101"; -- Argumento 3920 Funcion -0.26671276
  when "111101010001"=> s <="010111100000"; -- Argumento 3921 Funcion -0.26523403
  when "111101010010"=> s <="010111100011"; -- Argumento 3922 Funcion -0.26375468
  when "111101010011"=> s <="010111100110"; -- Argumento 3923 Funcion -0.26227471
  when "111101010100"=> s <="010111101001"; -- Argumento 3924 Funcion -0.26079412
  when "111101010101"=> s <="010111101100"; -- Argumento 3925 Funcion -0.25931292
  when "111101010110"=> s <="010111101111"; -- Argumento 3926 Funcion -0.25783110
  when "111101010111"=> s <="010111110010"; -- Argumento 3927 Funcion -0.25634868
  when "111101011000"=> s <="010111110110"; -- Argumento 3928 Funcion -0.25486566
  when "111101011001"=> s <="010111111001"; -- Argumento 3929 Funcion -0.25338204
  when "111101011010"=> s <="010111111100"; -- Argumento 3930 Funcion -0.25189782
  when "111101011011"=> s <="010111111111"; -- Argumento 3931 Funcion -0.25041301
  when "111101011100"=> s <="011000000010"; -- Argumento 3932 Funcion -0.24892761
  when "111101011101"=> s <="011000000101"; -- Argumento 3933 Funcion -0.24744162
  when "111101011110"=> s <="011000001000"; -- Argumento 3934 Funcion -0.24595505
  when "111101011111"=> s <="011000001011"; -- Argumento 3935 Funcion -0.24446790
  when "111101100000"=> s <="011000001110"; -- Argumento 3936 Funcion -0.24298018
  when "111101100001"=> s <="011000010001"; -- Argumento 3937 Funcion -0.24149189
  when "111101100010"=> s <="011000010100"; -- Argumento 3938 Funcion -0.24000302
  when "111101100011"=> s <="011000010111"; -- Argumento 3939 Funcion -0.23851359
  when "111101100100"=> s <="011000011010"; -- Argumento 3940 Funcion -0.23702361
  when "111101100101"=> s <="011000011101"; -- Argumento 3941 Funcion -0.23553306
  when "111101100110"=> s <="011000100000"; -- Argumento 3942 Funcion -0.23404196
  when "111101100111"=> s <="011000100011"; -- Argumento 3943 Funcion -0.23255031
  when "111101101000"=> s <="011000100110"; -- Argumento 3944 Funcion -0.23105811
  when "111101101001"=> s <="011000101001"; -- Argumento 3945 Funcion -0.22956537
  when "111101101010"=> s <="011000101100"; -- Argumento 3946 Funcion -0.22807208
  when "111101101011"=> s <="011000101111"; -- Argumento 3947 Funcion -0.22657826
  when "111101101100"=> s <="011000110011"; -- Argumento 3948 Funcion -0.22508391
  when "111101101101"=> s <="011000110110"; -- Argumento 3949 Funcion -0.22358903
  when "111101101110"=> s <="011000111001"; -- Argumento 3950 Funcion -0.22209362
  when "111101101111"=> s <="011000111100"; -- Argumento 3951 Funcion -0.22059769
  when "111101110000"=> s <="011000111111"; -- Argumento 3952 Funcion -0.21910124
  when "111101110001"=> s <="011001000010"; -- Argumento 3953 Funcion -0.21760427
  when "111101110010"=> s <="011001000101"; -- Argumento 3954 Funcion -0.21610680
  when "111101110011"=> s <="011001001000"; -- Argumento 3955 Funcion -0.21460881
  when "111101110100"=> s <="011001001011"; -- Argumento 3956 Funcion -0.21311032
  when "111101110101"=> s <="011001001110"; -- Argumento 3957 Funcion -0.21161133
  when "111101110110"=> s <="011001010001"; -- Argumento 3958 Funcion -0.21011184
  when "111101110111"=> s <="011001010100"; -- Argumento 3959 Funcion -0.20861185
  when "111101111000"=> s <="011001010111"; -- Argumento 3960 Funcion -0.20711138
  when "111101111001"=> s <="011001011010"; -- Argumento 3961 Funcion -0.20561041
  when "111101111010"=> s <="011001011101"; -- Argumento 3962 Funcion -0.20410897
  when "111101111011"=> s <="011001100001"; -- Argumento 3963 Funcion -0.20260704
  when "111101111100"=> s <="011001100100"; -- Argumento 3964 Funcion -0.20110463
  when "111101111101"=> s <="011001100111"; -- Argumento 3965 Funcion -0.19960176
  when "111101111110"=> s <="011001101010"; -- Argumento 3966 Funcion -0.19809841
  when "111101111111"=> s <="011001101101"; -- Argumento 3967 Funcion -0.19659460
  when "111110000000"=> s <="011001110000"; -- Argumento 3968 Funcion -0.19509032
  when "111110000001"=> s <="011001110011"; -- Argumento 3969 Funcion -0.19358559
  when "111110000010"=> s <="011001110110"; -- Argumento 3970 Funcion -0.19208040
  when "111110000011"=> s <="011001111001"; -- Argumento 3971 Funcion -0.19057475
  when "111110000100"=> s <="011001111100"; -- Argumento 3972 Funcion -0.18906866
  when "111110000101"=> s <="011001111111"; -- Argumento 3973 Funcion -0.18756213
  when "111110000110"=> s <="011010000010"; -- Argumento 3974 Funcion -0.18605515
  when "111110000111"=> s <="011010000110"; -- Argumento 3975 Funcion -0.18454774
  when "111110001000"=> s <="011010001001"; -- Argumento 3976 Funcion -0.18303989
  when "111110001001"=> s <="011010001100"; -- Argumento 3977 Funcion -0.18153161
  when "111110001010"=> s <="011010001111"; -- Argumento 3978 Funcion -0.18002290
  when "111110001011"=> s <="011010010010"; -- Argumento 3979 Funcion -0.17851377
  when "111110001100"=> s <="011010010101"; -- Argumento 3980 Funcion -0.17700422
  when "111110001101"=> s <="011010011000"; -- Argumento 3981 Funcion -0.17549425
  when "111110001110"=> s <="011010011011"; -- Argumento 3982 Funcion -0.17398387
  when "111110001111"=> s <="011010011110"; -- Argumento 3983 Funcion -0.17247308
  when "111110010000"=> s <="011010100001"; -- Argumento 3984 Funcion -0.17096189
  when "111110010001"=> s <="011010100100"; -- Argumento 3985 Funcion -0.16945029
  when "111110010010"=> s <="011010101000"; -- Argumento 3986 Funcion -0.16793829
  when "111110010011"=> s <="011010101011"; -- Argumento 3987 Funcion -0.16642590
  when "111110010100"=> s <="011010101110"; -- Argumento 3988 Funcion -0.16491312
  when "111110010101"=> s <="011010110001"; -- Argumento 3989 Funcion -0.16339995
  when "111110010110"=> s <="011010110100"; -- Argumento 3990 Funcion -0.16188639
  when "111110010111"=> s <="011010110111"; -- Argumento 3991 Funcion -0.16037246
  when "111110011000"=> s <="011010111010"; -- Argumento 3992 Funcion -0.15885814
  when "111110011001"=> s <="011010111101"; -- Argumento 3993 Funcion -0.15734346
  when "111110011010"=> s <="011011000000"; -- Argumento 3994 Funcion -0.15582840
  when "111110011011"=> s <="011011000011"; -- Argumento 3995 Funcion -0.15431297
  when "111110011100"=> s <="011011000111"; -- Argumento 3996 Funcion -0.15279719
  when "111110011101"=> s <="011011001010"; -- Argumento 3997 Funcion -0.15128104
  when "111110011110"=> s <="011011001101"; -- Argumento 3998 Funcion -0.14976453
  when "111110011111"=> s <="011011010000"; -- Argumento 3999 Funcion -0.14824768
  when "111110100000"=> s <="011011010011"; -- Argumento 4000 Funcion -0.14673047
  when "111110100001"=> s <="011011010110"; -- Argumento 4001 Funcion -0.14521292
  when "111110100010"=> s <="011011011001"; -- Argumento 4002 Funcion -0.14369503
  when "111110100011"=> s <="011011011100"; -- Argumento 4003 Funcion -0.14217680
  when "111110100100"=> s <="011011011111"; -- Argumento 4004 Funcion -0.14065824
  when "111110100101"=> s <="011011100011"; -- Argumento 4005 Funcion -0.13913934
  when "111110100110"=> s <="011011100110"; -- Argumento 4006 Funcion -0.13762012
  when "111110100111"=> s <="011011101001"; -- Argumento 4007 Funcion -0.13610058
  when "111110101000"=> s <="011011101100"; -- Argumento 4008 Funcion -0.13458071
  when "111110101001"=> s <="011011101111"; -- Argumento 4009 Funcion -0.13306053
  when "111110101010"=> s <="011011110010"; -- Argumento 4010 Funcion -0.13154003
  when "111110101011"=> s <="011011110101"; -- Argumento 4011 Funcion -0.13001922
  when "111110101100"=> s <="011011111000"; -- Argumento 4012 Funcion -0.12849811
  when "111110101101"=> s <="011011111011"; -- Argumento 4013 Funcion -0.12697670
  when "111110101110"=> s <="011011111111"; -- Argumento 4014 Funcion -0.12545498
  when "111110101111"=> s <="011100000010"; -- Argumento 4015 Funcion -0.12393298
  when "111110110000"=> s <="011100000101"; -- Argumento 4016 Funcion -0.12241068
  when "111110110001"=> s <="011100001000"; -- Argumento 4017 Funcion -0.12088809
  when "111110110010"=> s <="011100001011"; -- Argumento 4018 Funcion -0.11936521
  when "111110110011"=> s <="011100001110"; -- Argumento 4019 Funcion -0.11784206
  when "111110110100"=> s <="011100010001"; -- Argumento 4020 Funcion -0.11631863
  when "111110110101"=> s <="011100010100"; -- Argumento 4021 Funcion -0.11479493
  when "111110110110"=> s <="011100011000"; -- Argumento 4022 Funcion -0.11327095
  when "111110110111"=> s <="011100011011"; -- Argumento 4023 Funcion -0.11174671
  when "111110111000"=> s <="011100011110"; -- Argumento 4024 Funcion -0.11022221
  when "111110111001"=> s <="011100100001"; -- Argumento 4025 Funcion -0.10869744
  when "111110111010"=> s <="011100100100"; -- Argumento 4026 Funcion -0.10717242
  when "111110111011"=> s <="011100100111"; -- Argumento 4027 Funcion -0.10564715
  when "111110111100"=> s <="011100101010"; -- Argumento 4028 Funcion -0.10412163
  when "111110111101"=> s <="011100101101"; -- Argumento 4029 Funcion -0.10259587
  when "111110111110"=> s <="011100110001"; -- Argumento 4030 Funcion -0.10106986
  when "111110111111"=> s <="011100110100"; -- Argumento 4031 Funcion -0.09954362
  when "111111000000"=> s <="011100110111"; -- Argumento 4032 Funcion -0.09801714
  when "111111000001"=> s <="011100111010"; -- Argumento 4033 Funcion -0.09649043
  when "111111000010"=> s <="011100111101"; -- Argumento 4034 Funcion -0.09496350
  when "111111000011"=> s <="011101000000"; -- Argumento 4035 Funcion -0.09343634
  when "111111000100"=> s <="011101000011"; -- Argumento 4036 Funcion -0.09190896
  when "111111000101"=> s <="011101000110"; -- Argumento 4037 Funcion -0.09038136
  when "111111000110"=> s <="011101001010"; -- Argumento 4038 Funcion -0.08885355
  when "111111000111"=> s <="011101001101"; -- Argumento 4039 Funcion -0.08732554
  when "111111001000"=> s <="011101010000"; -- Argumento 4040 Funcion -0.08579731
  when "111111001001"=> s <="011101010011"; -- Argumento 4041 Funcion -0.08426889
  when "111111001010"=> s <="011101010110"; -- Argumento 4042 Funcion -0.08274026
  when "111111001011"=> s <="011101011001"; -- Argumento 4043 Funcion -0.08121145
  when "111111001100"=> s <="011101011100"; -- Argumento 4044 Funcion -0.07968244
  when "111111001101"=> s <="011101011111"; -- Argumento 4045 Funcion -0.07815324
  when "111111001110"=> s <="011101100011"; -- Argumento 4046 Funcion -0.07662386
  when "111111001111"=> s <="011101100110"; -- Argumento 4047 Funcion -0.07509430
  when "111111010000"=> s <="011101101001"; -- Argumento 4048 Funcion -0.07356456
  when "111111010001"=> s <="011101101100"; -- Argumento 4049 Funcion -0.07203465
  when "111111010010"=> s <="011101101111"; -- Argumento 4050 Funcion -0.07050457
  when "111111010011"=> s <="011101110010"; -- Argumento 4051 Funcion -0.06897433
  when "111111010100"=> s <="011101110101"; -- Argumento 4052 Funcion -0.06744392
  when "111111010101"=> s <="011101111001"; -- Argumento 4053 Funcion -0.06591335
  when "111111010110"=> s <="011101111100"; -- Argumento 4054 Funcion -0.06438263
  when "111111010111"=> s <="011101111111"; -- Argumento 4055 Funcion -0.06285176
  when "111111011000"=> s <="011110000010"; -- Argumento 4056 Funcion -0.06132074
  when "111111011001"=> s <="011110000101"; -- Argumento 4057 Funcion -0.05978957
  when "111111011010"=> s <="011110001000"; -- Argumento 4058 Funcion -0.05825826
  when "111111011011"=> s <="011110001011"; -- Argumento 4059 Funcion -0.05672682
  when "111111011100"=> s <="011110001110"; -- Argumento 4060 Funcion -0.05519524
  when "111111011101"=> s <="011110010010"; -- Argumento 4061 Funcion -0.05366354
  when "111111011110"=> s <="011110010101"; -- Argumento 4062 Funcion -0.05213170
  when "111111011111"=> s <="011110011000"; -- Argumento 4063 Funcion -0.05059975
  when "111111100000"=> s <="011110011011"; -- Argumento 4064 Funcion -0.04906767
  when "111111100001"=> s <="011110011110"; -- Argumento 4065 Funcion -0.04753548
  when "111111100010"=> s <="011110100001"; -- Argumento 4066 Funcion -0.04600318
  when "111111100011"=> s <="011110100100"; -- Argumento 4067 Funcion -0.04447077
  when "111111100100"=> s <="011110101000"; -- Argumento 4068 Funcion -0.04293826
  when "111111100101"=> s <="011110101011"; -- Argumento 4069 Funcion -0.04140564
  when "111111100110"=> s <="011110101110"; -- Argumento 4070 Funcion -0.03987293
  when "111111100111"=> s <="011110110001"; -- Argumento 4071 Funcion -0.03834012
  when "111111101000"=> s <="011110110100"; -- Argumento 4072 Funcion -0.03680722
  when "111111101001"=> s <="011110110111"; -- Argumento 4073 Funcion -0.03527424
  when "111111101010"=> s <="011110111010"; -- Argumento 4074 Funcion -0.03374117
  when "111111101011"=> s <="011110111110"; -- Argumento 4075 Funcion -0.03220803
  when "111111101100"=> s <="011111000001"; -- Argumento 4076 Funcion -0.03067480
  when "111111101101"=> s <="011111000100"; -- Argumento 4077 Funcion -0.02914151
  when "111111101110"=> s <="011111000111"; -- Argumento 4078 Funcion -0.02760815
  when "111111101111"=> s <="011111001010"; -- Argumento 4079 Funcion -0.02607472
  when "111111110000"=> s <="011111001101"; -- Argumento 4080 Funcion -0.02454123
  when "111111110001"=> s <="011111010000"; -- Argumento 4081 Funcion -0.02300768
  when "111111110010"=> s <="011111010100"; -- Argumento 4082 Funcion -0.02147408
  when "111111110011"=> s <="011111010111"; -- Argumento 4083 Funcion -0.01994043
  when "111111110100"=> s <="011111011010"; -- Argumento 4084 Funcion -0.01840673
  when "111111110101"=> s <="011111011101"; -- Argumento 4085 Funcion -0.01687299
  when "111111110110"=> s <="011111100000"; -- Argumento 4086 Funcion -0.01533921
  when "111111110111"=> s <="011111100011"; -- Argumento 4087 Funcion -0.01380539
  when "111111111000"=> s <="011111100110"; -- Argumento 4088 Funcion -0.01227154
  when "111111111001"=> s <="011111101010"; -- Argumento 4089 Funcion -0.01073766
  when "111111111010"=> s <="011111101101"; -- Argumento 4090 Funcion -0.00920375
  when "111111111011"=> s <="011111110000"; -- Argumento 4091 Funcion -0.00766983
  when "111111111100"=> s <="011111110011"; -- Argumento 4092 Funcion -0.00613588
  when "111111111101"=> s <="011111110110"; -- Argumento 4093 Funcion -0.00460193
  when "111111111110"=> s <="011111111001"; -- Argumento 4094 Funcion -0.00306796
  when "111111111111"=> s <="011111111100"; -- Argumento 4095 Funcion -0.00153398
  when others => null;
       end case;
    end process;
  end tabla;
