module decod_bcd_7seg_verilog (
	input [3:0]bcd,
  
	output reg [6:0]y);

  

	always @ (bcd)
    
	begin
      
		case (bcd)
        
			0	:	y=7'b0000001;//0
        
			1	:	y=7'b1001111;//1
        
			2	:	y=7'b0010010;//2
        
			3	:	y=7'b0000110;//3
        
			4	:	y=7'b1001100;//4
        
			5	:	y=7'b0100100;//5
        
			6	:	y=7'b0100000;//6
        
			7	:	y=7'b0001111;//7
        
			8	:	y=7'b0000000;//8
        
			9	:	y=7'b0001100;//9
        
			10	:	y=7'b0001000;//A
        
			11	:	y=7'b1100000;//B
        
			12	:	y=7'b0110001;//C
        
			13	:	y=7'b1000010;//D
        
			14	:	y=7'b0110000;//E
        
			15	:	y=7'b0111000;//F
      
	endcase

	
end
endmodule